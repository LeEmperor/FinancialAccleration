// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Jtf5nllPDvGVoe3cgvlLnNk29KFGQ8ogFOhA92RO0XGsXd7gqwcKDwY5cgxGiRfJO/x/N8HbxgWE
K/UrwifM6qva8Q6YMR1EzBhAqgqvMvjHNvqalu3VDyObvKFbjHLVIEppGACnovqFCear+4XjM/LL
q8o+dqKoL0k53UjDtR2EsaY7kvYDREgssxDRqumC+UYJNZwuixGu4A8AJ4hjLLYl86z57XdVHsiz
CBA5hnOt8s5GzyehC4WfnZPYk9Fony5sGnfYpwuXtqtc9k0vkSM7H7Pw8CQtNfpwbMEJTb9oG0yk
qygc86u1e5uFitjG605QztZBB7WTu6d4sH6q0w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
M+tMK2nsoSzMo32MyWQCve3KKM7ia4nbjaKn2tnb5ShThqPSlcEiP78IRxhX/w4ZtMnAkvn3pSsa
lRTiIJLjxQzfvPX0ijwc1iGhK9yjkB38b3x0j6upqvhUsnSJF/qnm5PBzSP2GrR4z2gRmIQfk8H+
+4Y7vetRHqBe3/E/i3w6J/s24dv6u6IFJVlgCjnxQPDQ61IYbuIl24ttLBtUdRV4oGOAhmWqGf5K
qiTTyvyFtLVMoa7blTvYzWLaLPNV+0lSgGcYQY6ct6bELHn8c4m8qbEsf2WzFPZ5DaEJB7oV4M2a
ZMumIk/UcKXeRbw/ZdhdZwAUNNWqh797XYJxGA4NDNkNhfQTuSvOxWPZKvxcLcMl+40MP4RADUzn
bM+SisywCxvBB9on+NpQl4SwUDcQVLyZ+YnNhRbRrvK0n1YRy2XBAHp7/ZAWZrP6BWGNfmd9TVI7
UWaQKyAFDwCa1blZ8x2SMU4OnngdjNmB7zuTkmQXnBKw+zuZGZd8Sw+/nUUTylwPlQKHw/gTXO5+
ZN12GlV3/xAUd+rmAkQvMKE4dsqQsljPN7DqG7YcckyTKIUNl6GpCnWT6FWPK4shBkv8gXxdQDeT
c2v+rCUHmJX53Vte6AFPHowBpCQuLZ6B4nQXB7f+zcDIb7Q1AFnHlibitBSYAsvgoFz4/iHeRc83
w6In/5v0q8deVyzeXGZcpYQje75uA7YkGuiPwfLcWoMxRCiMOEsjDGCj8dTN3xyhgg26dH7T/nsg
50z1q3LKeAvjgAgv2g4bzJi4hx5XyWg9cgfmCe/l45z8WRdpCcCaPzIO5qrFwSQdeHKUvi5cXRLT
09ZWPbAOeorZ6WOwFZ5RvUcvl9xVaBcJd6FXVJVsobA5ftomSXB8Z3+v7yG8JslucRZctQ4LuMkr
xpCylb9wMGidXkKK//t8M837rFsME8j0v9pZqEJiHBpO+Gxl4Ly9KWhAuyyRDsXesXNyHjPV3GnF
iQ+XGcWGWZ7JT7CUgvO6gDDaJfii0eUatKmc7fw6tXBtE8CuKNEAtEhom5gyv7ktRtl8LTxDqw2K
N+0XdUSbNxIGW0p+4V0BX9itD326zEYXbO4yMuNrhDhsdBlBJx0cjOvMmcqHQBNwepMhCOqfGXNx
C/OyK1Y2BsjpuUM6WzmtBg68NId7nsRRMhgs21Kynflp9yda5UGmZ9r2e8+Y2343KfP1/3XpVPV6
skC4kPLJ/dDgDvTH0a42iqDRY07B64PGQhmpDK1va8CCTbCQplkPrBcaylVHwoYgNPsK1xZLB8Bz
AwFXaSZ6c9pnTt2Nu9u6vX3wFW2A5C0uu9oHKYwE/NsgXal+nOSN+DroCwtgciTSjgX+QihYgS5M
/NDfKWa8UB8eq6hzZ3jS+4EJzX/D6tP8dVWly5Gtl4RMmZ7omAeG0qxtekdhDrSpKcywAW0Ap6yC
WZ9UwiY04QZaWxmQYnHDRt6oe+j80qVU+nM9f90m9+wAg2niC41BIz8TIzWVOTlp1gzNghDQXjAU
L7Xaveq3YDmYeakHnMpqkYPfXl4O1ZZKrNvFDqQiyhGYptMWBomslxVqISvFcEq+8rUs81HAyXKK
rZJmIXj7Ffpbv/f5Hrler5E9RfmCgntmLgmniqGXlBU5YvQu1p02YO1wdsTMgLDnbGUc9exQppQ3
GPLUgnCJABquOsE703FVwX3NO+JpyYWIWti+MlwBBqWkw1y/3Zqw/j7fXEcScZRg495M6fCJw5Xe
W/F95ZAEmPlacvKoQmzgQgVZU+QaIAg977CKj3v7XU2aqzcYntJKQR/0eqKxxh0naK7q7k6Lsudh
3tzmidDpJ5m9KyCflKsBPmfdiaffh/vdlHXlQWuaOUZ479K4hc7heUHqM0YF44rPTDeWjUeI5wFC
/ErU+150Nn/g529RPqpR9Fz+OYiRCf4OwDLKwbTMKF6uvyG7nVkdo0PtQrILCCDNXiNiYtIT6mB9
lktG1n8ilwP/aZX9z0t0WCNPsCPKVwizhuWKShXmHSxV+RZ+iSakoolJGYwYlv+bXdDrDrs63Bnr
37rS6fSJhzcAB6fR6mfOIPGsfGYJUWGrXUcPcErr4gRbipbyHNup3xlY/YSgpHTdOtuuPhK5djF6
DLr32kkAaG+G13NLPwYLqQmzImxEoJwnTDZkHl3lmaZSaK+FaHTMas2nH81tTfrEIIDUy5nFXSn8
yLpTXDGXiE9uxy+HVcmgk7GtcwJ3k/vKsFappT1F+7JvmD2GxSD2uE1P5MdJkEXSlbK7AlJPLO+U
RVgjoeqi4OzmHa+HdsT8+h0CHqy4bjdX5o8koFVQ+xb73ZLp/yxGllvGVziASolD4xerWkoOWqRy
hhqsAmkiHWNSY67xC9YQlkfJc8+QoIUvy4pmBgeEc3MQsCrWlePz3hC107e6M3iFWk5WODdJxeAO
nMqaepycE0nMf0G8JyPhARN8H1ZYlk1vZBzwAZ2lgNvUqPRavtk4yXdQ6fHTEEeDlR5xffNgoqqy
M9XxBtLn8art3ascumTgWnaZHoDhQMj2pwTSvezSB41NdVaRpryVqq6W8rnItyGEMoLefz4qh+BK
OlPfXBgmU/tsfrN+15w6fgdN2jrQILYG9CQViF4yelWzdjXkaBPkV9Z7/dxKR2hmgakdZOGzW/FL
rstSg8GuERka4qM6zH3xOEfIThslbtFLjCcUEkqOYXXRjJdlf7b02ceruorsydGadOwSBKDgUGrJ
5JoyIrduAwxE+yEXiFdZvJRcGxU8DacPUCeoZzDdQJ5X1TnSRJcDFLcLtSnFrXDTs2tLwcslC1hm
zZIu6eSiW2PLoFE6rOErGYaVHJ6aZpbe5BAHRbTpi+WOQS5GHslfuz6gKiogkLKy8gHi0UNhWXUH
TPYwpYB46yv+62dgm5cir8xvuPfjvRICaoM+LXEuc3lPV33jU3fTs4P82blu9h4Hb06Y1mJUJ3kz
6JdP+KVD1xYGpmBvPTg/VcM2QBkmy3F72ef/vhbWMIu/ynib9bmd3gXY7A5s7oM0khKcxrlgj+IC
Mq4Rk4Fcqkf+JUonE4uxIX0TJOp77lNgeGCgQPHg/mCbN+mXRX9k3qH4596+gF+xHiQ/dKmXCzOs
ugOORzo9WMOcQMBVI8BFF6ofPSJQKwBe3J6ZsVHskVSfKScT+9aZoooHOB3BgF7+49tIfHQyDNFo
IDeMG0Hmk9wwlazr+mSkIreID8if9H0mFqucpjo1patrkOEAZoc6r+f8myqwJEigLJy4GDIKZb0R
iRnr5HEQp1lJSIwiWnZOkGFyDpPGA+ZoZ5urGkKR2ntE2YspYOdmL8JjxbrfR5sAalQ3DxSTOirP
3zvBQsjS2T1MxEX4yPpalhUUs1hJnJVihFtu5LbYA+CfU2z+X9+dw7nNyzzRz3jUROUIfsOFrDx1
O9g+Jn1OThkwLYR1sJj3lsHVA2XDp7vpM0e/+mbV2EcBydY/nSRfozNs4v/o9KYa8js5v/LII1eh
2yV2DVssA05d5Gf3lrSLYgiYln2zyD3L/r9W/TVMQEWs1igb/WCzUt41Nc0AJcJK3t/isIKwOhbU
r6JN2rvMETTBfyBiZAtAhCZ/7QUDHzUw16jXe3URAlA5ZAeENobB/N1drL3OGvIaxoj3nk9PP8Gi
5PJK//R3rZ23n108R4t7YgyGFteODfU1/vp92MoqLyKGMQSVZiALA7VXwVQ5UWso3kwLxJM1Y+g7
PN2V+pLengGA4EGNyLiMMCcH21ThP8qQuBxdwZ1GJ7pJwYIXpbTIEnyd3dzcXU+LkyG9Z3sWFUxC
DliGL2lpfznfYNuiZkTNDxzwvVaN+7Rn6+aYmCygsO6bXhYZE8Oz5DdQiWBpqyBYFQinTCMai8Jv
9DS8t5EhzISqf0CeEzkRTE79Jij7faJOTS2rY4jXtsF/0xa4X+/Ck18eeNlhlVsp+NxplIkYvMX7
VovINZKE6TYwNr9+SaILly4WPOlqvH83fp4IlkmdRXJ7dpaVDGSs9bsg4HOxn9Kem3aPSz3emc+r
OffQL1UoDkNhOnx9wquNAcRowvdpziYvVmqBBANkn2isleqJ+k+WehKeJupKMrcL7jiJt5yJtB8A
6hQkV1GQ/OFcplpfMuZEGZUpbrGgU1Y53sgqHAMApSeKZS8zAM5/qQ9qILoFnXdKNm8K4aXWfer1
c5rYT7tppGzL86j5xfYfWzbshWOlEWFjAaZHd9T25O9y/NA4wkBbmunjROvzd1oMCFI8Ota6CymY
iXOPdprrKU9NWQhxmTJDgH6iWgF/2RknUb2oTbLj5BmQzIhNR83oc5/ZMrcYu2jPEQlzWgtrV+Gk
v9Geohsdh+bSO+61nkn+uiUSF6K+vq1VfhpXKiFCT+7qDvioJ6vtrp6cp588nyEbvxaQ97UsLD/Q
I+Ps1t6O7UtiPWx1V7muWaodnDtrA0RHnmDv6rJhcdj91NC+2MEv3x6Vv0uwyOTyyQPswn++VfU1
vi1CdRSVJ96Lg8gui7r2ofWaHZ6PJbok/+uxKcF+U02AZNB/tltkugG6kKX40hAPEt0m+6AqVkt3
hlmOZG/2W0u+UCR9qJE6M7GhuZeVN+lfcN6vs4ICjygUlKK3ahnQlgGQuvfWp1I7c+obzmOnt6ZM
QN8gQ+5EzN+zenpUFsCbKZsOyEVQ+MS/oC2BDR2KXjftGheBOQQm6o/ALxQfKZVECy1ru9KivCoX
EDkwrWP4m6AVDdEmqAYgOni+h4l4FMn+n9eUorDxj/zLjpaXws7vVRFgS+I2H8cmDvh+b7HiqsTl
aSPOcPtbtEkXL5T4BajUKoLPI19OJdbeIcHwQHZTBgVk7fGE/gTVak6ii22JasUq57Tgd905h8We
eSpoR1HuVuCkP0n7+fVE54OwW5d1rnuwmgn9ltowl7reVigiilBFX7Ja0ottDlaZk4/VOMa9+ZKM
XYsxV5yc7qbtpXIQTnH/kDYCVaR0DCulIAKEHJ2oq7yeUzvKIarup1fEQc5dAXW7Y1AEVh0VdE4E
f0wO8JN0QjjdpwPr20c5mmjeDEii/xaJsQAlx0dJUoySZ1XlpmJPnxT7T35hq169OoIKxB25nZ+6
EqsCQ/DcQsqXha+SwY4n2WfuR0ktp4YbCeTXwvjGCT80flOGsN1s2LL4vf+ImBeOAHsgj9KvuVY5
Ut088p7gsOxyTiGUoDPQXl/z0FpOU4R66SHqYqN8TYPji/9Nc0sEnDwRos+YusGNHr4LIJ274c7W
W5nTAPLUg67HWjQQwxrJo/PX6m4SejWMtPnIoNOyVe138+8Fp3nvhGskGi4eLjqwb2CXs8bGYcNK
wog5x8ppziYndN6e3sdTZkemRNuAnlrFwWoLEr3ozafmL4Gcb2KtFNaq2Fbwi0yowUt4iMLS2oF5
CwNyO5klS2VHgKIsR1S+XJoFcCxaVdxc7scoIIr0QIRQexH1Bfpxl+n+QUfkFV5DX1fpD+5SidX/
faDouf1aJ2zJVgZowoBczu0kyTfcuzyuleg5uxuKlyoetdgdhQ+XxWc2xd/MK25+D2v5qitrWY9q
2DjVlIb9awieONqYApFarliKo9SUTSt2DDR3mwmPgFl4T3xddPHCVVjsPt+52SkqKZhku8Ncw800
2fQpoOM7Wq/GZEP4UkJUWvZcx2pLydfm6tfnpVkpC4lI7yApxNVsp425aliVqHXssXC2i9imLoR1
Wdv5NQDHPWLGX0GCW0WYbeTvsQh58v2z2z9NVbcvNX6Z3rOJvuHngmVjweYPdUSVxuRJ14u/9Iiz
HkXBGglHawtkm+PIUdqaPACXVZwadq0FeH+AJ3Bjw507IN0n02ChBGMbUN/VWLIDAG6KPKVpHI06
j5boGNaizCyLcO+AD0RsU899lJ6MLWEc1cKRwGzHHr4RGXGlgZ3t1ODPxvENz+dVl8v+1cg1NXIk
EvcLePJtGCmM1BM+0qLBr1hL1kajgfu/cgOxlupf3HRLEZPtUZAPJwjBEF6hL3UktJSFVG/3KYTs
VczUNZwU65nlePvRldTpTS9A+vEVOWeG44S74xC6HTxQVNnJpOSvTnHgb1Be0y3Nm9xSvmiAqtdo
niwj+FVHefh+/rkf4RGQouwGsKlFyRixKIyAaZH+6tV6OrgCgBcl4zx8Z05n/OBM1COGk1oQCkKG
N3NNjc6PznDNJdyIUZbH9tjMs59rFUGgZURoX80MhYbN+9W5j6ZWBPfWr3TwC9gKSZi7yUaUq3US
M7gUQscD2T7VGq0aCVo8TOTb0+znpLcr11wkjIEaVy4+AKiIgjVaXjy07Rur+FKYiSvOCiNhNMUC
/boRvd1G0WcFNHuqPxdnnF1VjtQIQhyzn4u9mUWjsgag9ILMz60ZFXKponPuLur3spPOW8tzUJMP
Cr2qvbks+d0T34V8o1IHVkbqsiJXZxLDUCe4XaJLnyvKrYuxptfRlI4cX4Nx16sayYw3xy0oJTZf
ppMCKcWC79lMB+R0ZN3qwEMTnb2BMb9++SOWo8B5UhbB7jfP4bwHp7yz+OApsQdsbvDdH5ZrSXaM
2TlUtT4PJF70qmXwepPd0aG/KfB8dJIJ/YjJIqUgA3Vq2sJZdrxShtoaI3GfxdY7Vf9nWW3kcpjg
9z1rXi7j2s6X9e+AzOCSIjb1cg/6QBo7xP32d+ImrEn/tBu0csII1x01jRa0NfJ4LRg/qPwyS+Ur
3vSxbCdeS2Ob2UCLLt07TI3NulTtywjdbewIWhGgwkIuhGNL72kKbkkSZIiyYtpLtiysJYaTPA8f
XsFbhppVUvVBn5YWCzaMxPbjrWqbcp1u478Do94OhovMCSWP+yI7+q/pslGX4+2Y4aXATSrPcHY2
70fa5dSlyXMjvbAN5D0VfYYoUW9bGwwYZ8GVepXEp9ppxa7DnceXqpsFD5NW2BBsWKi6C+mxSaD0
TP4cDwaFNfhAQJTesOHBVeeCYh1gc3aQFz4nGr8iuxoyrctUxvew11bVa86xBGfZ6TUBKYviFBHd
lDXVX5lxcYVwE4A4byQYY02TzfMimqSYwcecio0uu/kxe3JFWd1r2rl3tvQQzNoxecUDIeriYj3h
FNwDdwiUjd2nYavYAYY0sw259/cOvV3i+gNHUpQOW3e6NCPpU+YKfxre8CnWAH9c9rmDJyue3jeT
pmaIDdCQwROy62SqPedoao6O6Si2Z6ZcoJ688Q0SswzGmEb87CxJjjmZaVg5kYlnWbouJfRehacQ
sOCZ1C1Q5MvJbxMtmaVdaW/WkZR7enmzO86ZCjV/cTOfnPjEpX9K/BGFMmATRTJkBOAOMb/JO/rC
r1EKFYOzCAFF7wI1eVySl2Hpds9xPwncJlbXCWMAxJCVtYY8TX88ObzIXWaMcu3FO6+M0KGjurUp
saq55QL6izAmz4u9zvlfhCjgn3XdroGM5EHtrnsIjBmMJNjguWMSiKKi6lQJUv10zZNlFvX5/3/o
hglsp3WU1uBcsRBiii+Sm1PP7t0xdNMjv/aEMekGKPh8Zx0LRzBPa2bmnq/g5l25eQ91hmWP5nBn
Gff5dL/StTajMXkach2Uw/qbqdbYe9ap3tAlS1gl6SVq3T9aw2ocUCNQ4kR31wtSeuKb4BiQ7NBC
R1LTp3T0QRl2WC7030uM5SNUcn89YDwoSUc50e94jpOMk90Be4VeLm/i3x08PFPfU3gKkqde+1DX
yxg6
`pragma protect end_protected
