��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��x���9eS� ]�_g�Xh3��1��63�A�1{Վ�eb��9��d8_��g�G�oWs$㩕�䫀�*Q���7е?-�@�Z��.޷�0�Ȭ�*
XL�1���-ec��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^�ُ�VT�T�Ov�k�UzI�n<�\�-�(�6��F�����UP�3`3��݁����T�+`����nӗ����
�-�ԓ�?m��`���t����ʀ���K6#���F���e�zlrћư�r���Tv�G]��s�hMR�}�`��4 Uv!ՠ3q�f,E
ZV�e���#���L#Ŀw��C�wT*=C�ʋ�ȣ��# �Mc��^�*���ra,/�fh@C�/��R"w�YM�t�� �#���_z�E~R2u�������	�y���K+���xXzmp�ҿ-�

L�Y�)���&2~0\�]
�Ij+�.�����~gC^F����P��?L����d�����%P�c]	
�7�u8Y��i�$�M�Ɠ'��Qd;����6N�U	�9.�5̜qp��O��mt9���#�p�-�)q��o��,��)b� "����x�x�NS�mW$b#:a6���]E��}�2��H��]VjP���ܘ]>:~���]��<�!d����ݱ+����t���,
���3��v��M���o�"5�X�:�����J��5���"�� f�p-���{2�_��4�x�=�I�E�����8Pr��P�'2��R����A(��z�b�T�����&�l�����09��hyl��z̾!���{~�;�U_D�.i�;�#2(�&L�N&*:��	�P/��@
-�Ҍ�Y��?�����m�7*�z��U+��u��`�s( ՛I�}��ߐy�L?m����!���]L��SH��7
e�v��eX��Cǚ9��K�h��/�Y&#�~��cth�n��E0��0�[�����<i� �|�|���,�/���@j����K�V�>�j�b{���M���B�˕>ehAX���.!q;h+ǔh�!��Lg�,)��td>H>7"�nd�vmzj�h)��!��pK� �x�8�\q�N�@.�8!2{e��h��֣�>6=��G�4˫�L�=�2X��&5������M�n۝���O���7h;�L���TÈY�ӧHh��'2Y�l�l(��z�����t�d�{����4 ץOxO����#���Q�7'���S�%��Ih��ί<���Gɗx�N�{��0�BS�w��+^p���Ձ�3r�V�ZQ;a�t�Fk�b�����R;�S��b�p�%�]�2����wa�f�:���}����1��=S��~�T�����I�E(g(�D�o�(ޏk�ud��8��!PBy���F�&R}#��1�	lՑsl}���ZQd�6[
p�B�UոW��8�+.�1��,��E�gT��wč��,�T�B`����R�H7��G��b� �h��������9�sj��g��O�d3sx�7��3��:D4�pC	8�����Ms��7N��r�'���6��6"O�ZJ��0�b]B�G"�W��-V̄�I&�[��nm�#/��Zm�/(p�q��X����BC*���y��j�f2^Ae�Q�4\�ʇ9c��iiZl��aWw�MX+�+��0��?�?����!�B2�G�R)�XQemD)��Z��,XMai�2��>���mO�D�n�٩4��R|�yi�~�@G��^v��ƒT[���#�{��:I�Ls��l�Y�(J!L>��9�3o��e;�X �~ L�r#�������i�a�]1*�`�8�ê2��:}��p�{'���"ؓ��U?�!�!3^��	�Z`��������=���F��b��#��}��r�xf�	�C������-�]s����Ńʹ����D��@�.�yW
���&�/eJ�Cf���'?�HF��o��(��d�j�M���
���`�)�6W������:Χ"�GJ��[��b�/�{�.�Uz�(�5�cp�O��3���r�t�|��8�(�iӐg�?OsnIa.fR���8�n؏,y-j��֭�'�7k[�$��>�u�_��z��\)~^��W�����#��ǅ����Ɓo	�'�m�	W��i�D�0�In�;m����$��ǿ��Ti�W��4�x�V9M+��9ߑ�Yԁ<*_���{��7��J�VD�,mDբM1�0�P��^1NY�I�(�ծ��OY@��8Ao�-���1��sh��������'����S���C��Ӛ�+@���FO	�:�>�P,������fK���KV�����E��'��b��t�W9}�]�.��j��F��,���+��;�vӖ�ISF�cR�ZFks��������c���vV��A�g�L^nZ��yT�_�#��w�Gv������(��YH(~�v�64���z:H�>o��~����E@P`��b�/�H��}����uS�2�N��S�u�l��s��y�R|=p�)�N@`�\!��cV"�wRʒԧ����`��_w@3�eR�2�%=��R`�)�U �⯉:|��4�<���WX��7�c{��)E�i��V�����e�q��8*ϣg��1q�*���H^�8MbP`�,�s�<����NW�Ťw���e	9�I�'�X��Ԕ��a{�i_����丞?��L�Y.�1�$���|#9�]fr`�x�����E�D��	���#l�-J� +@x���̸��}�7��.�ഄ_A��=��][�zx�����Ŏ6|�.,����/C��K��6�!'���8i;����zz���^�� �Vt��A�u������u����р��Rg
:��#a�G<�� �G�f�H��@H��1g&�r�i&����L.Mcw����c��I���@8��@�!�Y�q�t�v���WoF� fS�˹�L�*�ù���-��Qٺpu��T���?��.1+�aW]wS���TСC�C빺�6��6����7!݇[��:��T�8�ڕ��R�)>�gQ11��}e�gU�#<f��v4����e͒i6HԹ ȋl��mȶ�_bP�����67���k!@�ց��Jo�u���0
�WS#{
�]�@�4�H�jS�@���t�d��ԟ��4��G>��V�j�bR�
�)��e;�wc\���3v�9̈́ZQD	p��`�
ݶz�k��J���}D,�㩣x�"���U����I�aѴ���%��W����UP�p�� _;����!3�sO�|8��\R�i��M�c,�}H�����G�'��TQ1F�� �bx٥�`�x�0�b��sF�G!���_s�q����<���Þ/t�'چ��:��|�4Y<���^���j���M?� kRl|*>HLV�{ �)ʨ�T�4�W�����>][���g�O?򪫢���F�$૘g�|'��R<�L^�Z+bCp�|`��t���׊����D�z4��m���+;�	
jw8�q��b�z�BO�zͻ�H�,�m<�Ec�������(b�W�1羙��$�X�|O���G&k2�
�YE;�����G�	V����,8e�ۣP�izT�
����0��JE����ͬg�ێVN�LL7����X��^	Q%!�;��(�\/�����|B�\���|e3�����SP�Q�c�"ASK����hJ�as�)Yb�]4�n�-&r�ɶ5��\M�j-q'azj�ĎNU;�D��3m���_߃���1��o������N}��-��v�k/M�����ZQ��Oa!�hF��a*��Ȋ=O��~t���宲�C�����Fp��3?��]�a4VL�9��n�L�%�[��%�ԊV��2A�2��ܨ��Nf���ߡ�'B(�S�3�
�������R�
�z��li �1Ɲ�P: Cm���{��z�XF�&��ϒ�^��ruda\"Yd��Լۢ?+����@߭��4_���L� �^!f�S���5఻� s�~�_(���Qke�nY�}5{<�����#T������ݨu#�Ð��KziRë��y���\s�V܇���[��߉o� ؊�����i�U�J/�d�H�P����7�}���~Q�KI���y&,":�ߪ�����(	��D�sQ06��-�V)[�l):\�V�`RX��W���&�XJ�U,�!p�����"
�������˟�<�k?@�O.:#�3��ti^hԓ�d5�xOs��;��7̄���J����KR�:���@��t�I;8�������)G�[)2Ү�Ζi��x���#W̅,�3�LN����S���ov��yvG8�;��ӷ`��ߞ��r�` ����܌��h\-wH�e#At`c�6�$~�s$2қ@�2���G�,"�0^�3�3���7�y<2�}FX�rs��41c�sT'���T�>���}�^�L0�}�a5��'�fU�U��]e�1����o�q�Y/�,�,_�b��zoY��zī��}���2�ƪ�ު�����\P׬Uα�`��;]v������Ya)�Y�(;gi������?G��\?3[����!�r�U�6����N�9}`��u��dV�`�v������j�`�#�ȧ�ξc��t�WY�CY5�%Бۢ����S��r5Rrm2���˶�a�8Xt�xu&c#]�����Uda0�0$��V��pR��Y���U�Ռ���Y⤻綈�a�i�㷚��'��bfk3f	A�I���L�*�F�G$"d���7�����ruI�s���[M�wG�i,����!ԯ�z��m3]�]G��ꎍ������i�m