// Bohdan Purtell
// University of Florida
// Test for Board

module test1 (
  input logic a,
  input logic b,
  output logic c
);

assign c = a && b;

endmodule

