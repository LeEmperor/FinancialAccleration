// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:09:49 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mgd9MS1bhoumixKPQMz4d/zqOOUYCZBIuGJXy7D1WD+NlL2SwmTsfjP/xRj6n5RC
00RUBptCMU/CwbVjL9YMAVYyVAweufwlQd6xzWAcSSmE9D7qk0ss1AilPXIBdBwR
FVWr5GaRN4NHhppGdHPjAx1Js7iLOM1CBRz9/PU5/6E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
ZunFjyuQgZB/QYPt2JawfL1U+LcI82onROanDzaKZpOQ4CBVr5XK5P2xENjwKRXo
O81kQXOp6QKHFydDBMYrP40/1q2rBVq352sl5Pzin4OiPfcdn/mI5iDooZqjbUjz
zE4y7Xn9+aKyrX8DiO2E/WahP5nwYQvjzdKNVsgUavboSA9G0opsgL/HTntMg9EZ
2Zu3Yb9tVD7o1RIibYcXZZ7qZcHqezfSPPdfkHLBV+2mskQXerGkbG0V8VN38yqY
SHizvxkBx2m6gMngB6GZsshgXFX4T8PWhhjoCFTiKMte0GBd7VbA9mn5Y7TkQjq7
i4SDIHFCa05vYwWMi3aKrJKZ3RNi+vCnPS5G7Vo3smsubvp+zLCq+4FmcBkORCA5
mCUdGd1KFsx0oH9fGs8Dvp/KRgTwukteICpCBzxlokzLfQvBO64CMxph64c5BqzD
PL7xPcOnRtB0/RrdyeD3gl7MtkEAaboMEfWcS4N2Jq0MfCV0o0safN3KAvyZZ2EW
nWPTF+QnY8wmurHiH+Mr9tGvvN2A6xCZu2Wk6xPtOAcmc4i2IUfON61B30VOdTWz
+Ea0yFhQAZxnwfvSzfB70YWwjsDibfHDnRONPECRgxDHLG/Agtmoy0MERqWq30sS
kx4VEYM+ld2JkviL23t0lSF/JjQmmeV83AGrAY+g1htpBDopXfN3eD1RaPEzmaOd
uELktwItHacpHtFVaLfecIqTByI0RVmLVZhQ0lrovgUKBSJE63vNxJD11ffZRFJM
ijqOLpKOMsR/nqHmS9Ie9CNsC8sDPXNb78P+yANQzQo2S7kMOo5bcQ5tut71YmXC
v+7CW29zgRNwSKqXrj5IJvE0qY2TWOuLLY4KqhgIZsI0TeN8X2zzxh/U6C4kwwij
nU3+21IolXY8BLNXoZ6YaYS1lIYxnPsYvrvt6lCoUYQUuxvQqTdqgUws025UaXFb
R3rfvhin+ks4NmSb1jfkExd1H9UEY2TGnZKmzHyo2JVVmtHLcB5UwH/SckXCw1T4
1AwbbUhfy3nuvKWz7R/JtAZDv2c/J/D8LBJNnj2ES0K2yLYTT279gPvPKKr9jkff
e3hrptsGRbE/6J1vKPRyfhnCS8/jVx2D2PEidVIWhQ2LNjLM4kb0Am4W+9r1yG6y
FM0RDmh7VzTf4r9FP9+c7rWs/Bslds8M6WPa6HRlh3N/Khr9ngKnJv7S57ZRkReL
8veGOGeSQSnYdD+/DfB+NRsZTam5xTtuJMotn5efogmKhBEEey3Q7zkOotavrNpQ
Frq2n+jljNRm64MBCaQN09Q/FRk1i4sZ6eOJL0r2ntN4NlT39fh0wXv8ghPOaI0J
23k2Suir3OsA4+TFf6ZCbfACM7nAjojAvdWRFror4WWj+q/1VLKVE06Hvpg/Qca0
++3uyJ4/ZUptEeIIUUdhTkfrqWnzt5HrMb665oCewndV72AdJd2s9pIjbplna8dk
sqIEyLZ/HOQmZCGGtQkfczsG5GbGpIpp6iF/5tidTKglTJRVCiYFLQAgBpYz6MNv
ChL+WGK2IUZqPZ9XVb66zLlifqs46PfHVWV7lUCviUlHrKZVteHQPjBBMaIkvda/
e+Zs4xrJT/MEMQVcnuRK7CpETGmBf/llKeJpvLZTEmbGA10VfxTYckiB0zxLjDtS
Goi1EmoQGaBGoPsl5jMwoF6U5uQJCtQFcykYBqfX244DjrSYNN6563j7EiuXRnVI
imvAJrC6QBBUfgqSgKUaHvaa7GoZ8EorgLwL1Qdaj5Ie/0PvMmdBIGKox3Nj2DOP
rT+WiplEYspdj09KuRaxrDXd3Abz0L4+9xJaI/2xkoSTysDfiqI/FFJrnTNk4kad
u8J5Jwxggi/e+np8lz7uSWdI4LtICFv6IIOrXG+g7hJTechkgzBFGFucEAzpewgB
x/QTbeDdnwWROA9l5JLGFYMtE6VFCrBTwdgKTd6ZgEWM8Ol6aAyoxYiawU+IuIo1
/QDHXr+Y4+iHcfduftc/JTPGwEzrjX0PjshpGAMeodc6tH+anVkD9crJp136xmKM
letsqIQFQF/btx4WxDsHe/rv7I6dBH9Ph+dSg39vkU/N7rvgA0eBHSwF1Hp1IKGF
czGA0Yii99FqiEOF7XYmD/ENYAhYgTD5v9Yoh2hoFha31dnin5BiOSxXpBjJcrK3
TE0mg4hgH6XkLFYNx0mUDUlfCUheq8uwDl2HdPiyUsNwtwrD+UDg5yAudk4nl9wb
qboHXxs1ygwE6VUaYdTl5sY06kwK/uhIOFYOh3erWfjf6fZs9cr71v/OSMSR0PfU
EqyjKwgRyHg4DJhyjM7hkvDAArBTn9QhjQJHa+ub5QAuR2+/tY9ZxKkN/AU5g4h0
s9g9s6kVzdImgi/MI/8U428dTAvW46Dlu9JeGTDN0VD9NrTwIIpSMZdg11Af4UA+
JfDNnHJVi/1T5S6jDckHDkZKuRrHxSW4rRY7rQl3mT+pkCabDuIj4C1GcCE2o0Pp
eBMuf/YY3f1pMx5XIC/IbfvNWNVE65WOYhEjRbzNeLjznt2XM2zPwdgCjMnbHgJr
sEriknbqyuwDSYAXP/LYPhGWOtDnmSiFhgAIOcN7mLXcENxg61RmMPaTZL5fc7dV
R8p7ZRbQEd5DxcPgst+I4KMrqe10rwNr3g9qbufreYNcISLjxQCt6mlyR9zA5csl
r8V4BUcaEvN7ucg/hB71Anz0hsW6OqIbcEUiXV0Hsn4wZxAbArRc0q7FvhGPGl2b
YK0uUSuUW17W4lL1R8vouuF7MNxH9yRUOABt2v3O0kXV+SQW9IQAox7JyPKK06WY
TnfxYv4UcQkkY8yCn05sLzM1zBltWLyIZx437aTlX+0GlWnOglnqnpsng2x5ynot
5LQPTAt2X1nAPTaOdBD2QnhneGAbXWqQqkY3NBkaPLfZph5D6vv+H4aPmvZdvSFs
8zrXsD+zxIpf94QHNPthLmtpTI+hB2nH3m2k1JLfTIoVfuXGDdJYavXhsMcFMdxL
48gTIMhiN8JzGp1G6xCEHxEKvGE/MpCpgsipR6o12yQibYj4z3u+O1DNVpnrM8Ex
T/j8k6lPAQ7cu6DplxzgiwGLL+8yd5uaKyPO2mrKKhn8VEhiFaW2TA9BT30SswzP
dZ9Uoqun4R9AmHVH3ApKZvkYA5WNTyLCPoi16xdekvBgZhrGqhah7uBDaboSY/ID
caxpDUu46KL+yqCUv2YS1u+mxxrSnmXbBEVNxl7w2VXhdNjav/F44svwKfvw/lUj
Vhrh/9cjUjcNEG1agANInubKeYMZdbmdMJJN89Or8NaVxWCKS56vnRwlRgXWNixK
FisOydlHY0L8diSQt3dg6TDpu3P19UgPunbnzSCRthZCbVFLPS9YuR48ELdWa9kG
QCWDniAv/3qRTb0pk6l7OFYeHMRUAKMF5MGFF3rwz9ukCacP1RsI6Nc6e6OjPFaH
qVYGRPPdbUWbqtnQsLN5macr3WpcfboAutrt0GYWfAYK1rqcZZfeBPECmRoPF3v9
zeZpb6lxyUt7Qqv1KLbogkanpUbV4sjH4ZcWCVC4Mu9Ood3TZFyJSh+Fy9ZYzOIw
nyObTVhDUdPxsDVeVbdYZi62hyrelcJf19siHFQY5+ceDpssPmU+Mss/C+93FZ+e
ls0bXRpUOFLuKN9b3xixVD5urY6FzI3GGTLqvMEMdRwlNSZLcHmGYWiWgK94txNf
Vamd9jrIE63khH8acw+aDcUqtECDqZlY0Nhbfg0VuuYPL4H2RZzTJlJ+YAHgoOaH
PsAtqQ5ywknMp9Ki+/1Ej9EkeodfG7H1FIESqV2OrtQrPc/MeW7SBG+nCzqsPKpV
kzGQyPWJrDf3Uoa3nPisv/6TNcFJWxSwQEmi+MLogm9A/RS6FnmpUTbnbmHEIO70
JwRKY5h2kq1EpmVL9RYNlwdv85kaodRsdmTJ7i3SM2yT8Td6szgm7HQ09UQNXpYW
pOYT+2GdsFJy9sKyiT8t+hFL19xq5e4TJ7+OFTsh2SJN0xOgZlnxOFw2Uebp3Z5F
2r1sQRafCIGWEMNlRsoIjcozMzdnOsjx6wY8fZwlM6tnTO4PE1RoGrlfjJDDYhT/
5o+H1WBuia/sDRGLeC2UisIUk3SDbQz8f5GBmJh9LMqtD5XV4JrE5T9GriIlHlpN
xd8GzHJTXuMVEYmh1Yl8gHaMjgmYsIFW3LOXhG43gvSbFBIdrGTlDSL9L+gd1d9x
i8bxrrfKzO24/NqSFfgKkYxEirEf2q36ffbfZExn2TxDhwMdFrl8EXrdRaWDRXW7
bh6KuXlLvApDZL8C1EeVQO2VFa29AWDkpXOXarKUjf/pCMNUAX9zCna4PMMGb/n1
ZEFVDs1gUeej6LYKGafVjbSD4fhRiL2kqB2dQ2nbPiRUG6+MY37nbLjeoPxXDWtV
JU5mSRi1ntqS35ftb6DBYLoPTfz+0rNxl4FT8h+9iavfa4d0e98kuCKADTiyUpaD
rDqNErqcIP+Q9kvAHtahkB5LoW1OyaHESVScHVKWI+qMKol0UtToL8ncZtO7zJPX
bzpbZLAMCJHSuaxVRtGW4+GSbVbDaHIXR61srTWdYkWt7BWmjnfsgBNbj6dGTie8
4mEnetrmO396al7NgGHAdyEPxPZSxXi9P6IgHrFCdt1ikJm/1QuPmTBy4AiLQA2O
Y+LOKQYQZ+Rcdmm7JUPSsbQA7dO0+tbcpegMqztCNowrtni+Mln14eRwNGDLR/Qy
5qXiTFOxAm7jZl9JSpLmFrbcfp27pcdRotP7amDGnqLb3eCm0TZp11J/78IURJGj
RHVqnW8+LPCpRGkCsn+oQcAkpHLPcFLalC5mCtqQ2vqDrGS8pB6QBtIHgncq6pDv
d6m9KuyYKt+46liTLka64ZbcAi5cQ7c3N/6TRwu78cK9P3Ib2k8kgbxF3nmP9u/F
zL8Rx/N/JLWDRfivsEupv+NnbBeAQuxQr1nuFKt1CyZ+tSUDNyX+1h/NnBcuAXs4
gu3zJuvCpX/q6auqcQEwzCAW6/koRvjyFYlTbh3DaAztpjX8EiJzwGTL2oDmx7+w
I/EA10BNWzFN4PUmWbRJA11Z+pMcdmWwU00pPUmN2tU2ftIGwKQ7IEDDeIDSIzHe
bMe0Km1+U9siumw+WbDIJ0EM+bkuyNPoEZlw0l9+JWPTlP3mV19zJeaIYZgiweoC
H9hqpiaGcIKIcW/mHsYQgNTj4ZiV9Ypcwq78OiBX8TDD7nmiQSGB9KuLNfVUcKr6
w2UCiglVLBWOw4yxzODebWDbY+/O5kZspEkAoeH9PDrE1NqMOdhqrntitduhZQ18
pS++zmaVTO5MJMb9vF5Owh1OTxR6GBF0YJKtadSMWqNYiFNSf19h9O/GViZ5kZS8
zBzPIFo8Kwe5mEzmxC7X6cLctsPKpzu7d9tjASSz+VqtblIKGRlwLd6QUUe2s0CO
mLii0oZ9c8Bf66HEO8thkaIgDo0CKzqyZ/CTHzzNNLvXQVhTK6QL2Rgeo9TYg9Qf
+8eHd3hxL1Re/Qgdhn2USRMCR3NM/DgH/XR2mNJuuTuRjQPaxQMRC2D8nr0htlAi
XtfLQ/6aLiQIGu0WhaByi75OkH/IqBzp4lQJdKP84eFIMdqtlKJquVuEvizEHb19
etv+E4mXz1OYxHEisvq1B4K0f3kv77mv3OITvyBMqx/FBlOusop9gtVdtQyMclpo
4ApJs0t+QxuDiimqVkQ2Up5rOsC7utcFgm1brp1JPEOJuZq3MREsnWhIgQ+NZbyZ
Y8miNZFd8lXQzvQM5xstf2P6z3Wa3RJpXUKcsBHWF5r003FynaRCvvEqP+CrYFsK
DGwus6Q7UTB4AMGxAZJnNwtwqRAzB4u3mxFXQkY/Et497PzlR2i7dsg8Z1Eir/99
mOWA2TNa+fcDxortFdtRX6BTNFWqHuXQQeRlAutf90+dH2eyGQlTwZPpXAtraASS
r+5gWOPAOX0Lhdt7p27ev7o1ETVbd4GITgnWXoZKAtOoRPj3tf+fPbvtEOqWnKG2
guTP0M6iszOUHlxOHkYAoxsqaDAB/5Cs7xONggVV73mzZbgfqtRnL+xLaMwqH6W3
6Y27h456J07ud7NdsUI4uweWgeodt7d+NKJ0GDm/o3hpuycTT53xmHB74AWAFhu5
mjzo5cY6vDC9FnlotjqE1XNpRtfde6of9xNQQUuuQHT/HxyGU0hYd/ENlErNlrMV
GG80Gb1QNWC/fViBPJOrYRSG3Tjt0ldRKOK+uYTVth9aqXZnNGNAklAaQnwuClcS
f/g5JxCQhzOCcG/9gi2WJjTvjk+ky8tbMtMehK5s++4+s4+ra1/aGSwP/1RqC4w/
oIbzuXhSSz4jhPDt6P0IKB5C2zsWd4g4p+8E8eaynxn0Ja6NezLcOC8lIlX6tHHX
ZtPtJ2KV7ITlAwo+nu3OzRlcm3mBm9oSzBtRqVSIXI3CN/BPWzL3b3R/lrKiCGUF
mwyhkSB6JPed23mko8VXSkENPYSUF2PBVFbEogf7C3YmQuHWcyyGomYrNB/Bn7Lj
deyVl/mjglYGxSP8bDq7yKpDM0DxVIYTme8RIHwYjlRx0Lx1F1xemSGX30SgqjvV
VFkz30BtKLXR+69qfjjWpBvePj2dTj5CiDaPKHt0WyZ9eSvlGQXctCqBrZ3fmVyv
e7nNUxzsKWO9dR+6J0/JSU7MDl0tFKLBZijohN1yXnE59LIsCGD8IOqiiNp6CGof
0Y1eK4YnKOetB2EZbtcFTTDbWvttA4RcEU+RpDqEJemJQNldM3bQt7MhUHG2rsmn
5Vf1QT8ms12uU5P9yT969KIJyZZtaK5N3LAir7mZWC6Sl7Igq3I6NRji5V1Ajf7s
iq3noJMKXdnY+eLk2U2U7dZlbfLBKOkCSigvSsWYE0RvCnRIXTheffOC30/AxajA
OorL9QjR04AkJrMVZCggW3ZiW2HyBkJMmDQn34cRU9wHEkZ+r01i+Nz9hqdEMp5E
owWaq7JdjvACx6h05bACuEH9eoFxLQO+tgxlTlqWbrbyGBbjAT38fRLRwR09RwdA
eXb9IHkrrjBzPSONWXBcgdrG0Ir8k8IptoRGjSkB+dwt90DrobiXoCIflZyQtH2c
zi+TSKXVbxLeM8lgOQmn5g==
`pragma protect end_protected
