// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
jU6RuMrNyh1eIwFa+uVCPgpTPaEDuNek7jhmOGxuvMWv0g3jj9h9dwIZ9YSVttD2/nEHBgBCQsia
VKDRaS8q45KmbaVOeoJz3l4VaBA7BEw6NXW+PIU4nWlBTp+KZ09a+HXSBdIviFkLdowOHpLyWu69
Psm2YkkG2LKD22B7FfhuAzyP7qtu7ajbr/BzxQy9AvfNig0yJPBpyUW8oZaEJf9nASgrSSG8tOns
h5RLUui9y6Srss9TGyMu34pVP99jWrRmFG7Ldac21dAfnFqIp0euu+pPJnh9sPC8vQ+RLiHjgpM4
t23qwdGwTI/IcVxsQWaWHmt8Hb8jXn35+Mt1yg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
JLRJvhcytSV0PTPQokMGs227GkvpVdSU7Lzd1N6gGpDKmgtjiBxCkhY3nFF4ImsoHJUig1f1FIWf
RnYUwN0YrwcnZjhwUY+60J979qWJklbnJb42ol9BPlfrp3jkMjIqZgV1hZTct9CjIB6KlzVMEkX1
Nrxm/lh91932u7ORPq72loWqrLxZcIDiSTkto2IZ/r9pWYj1zsaVAT0LlLDNGadqwoGss1gs7fAc
kzLHwQXmQwCPByvxTBnKHgbm5uPIh/EP7JnS6GYw0MsZCXL1smUMdyzX/QC2pKKUFBa2vxuT5Xa4
eut6/EpQO+BQ/0JgiVk0fxmaHaCydQ09Gm7lIAKsr6TgUhHqBizxVuMWxWjDuyffh6asD8Ka53DX
8jfy2KDk1XQpxyEYrcxj0Ne9KQPm6nz796sdeM5KR1E5RJYBxMh9OdSnfALgk5O8DZMPR3gF300V
nFQqHw/QlMsCoO9qo+d3YcocQzlJIPDJ/48sVfzvDLxsfWcOk80f+fcOowDdpKI9hIjcicN6qLHK
b2N8pbK2C+PZxaaH69pm2D36xCrYc4d7Jwu7tJGyCVq6j7h34JEz8We29rQznqH4goqahmqZjfqS
8G01+T17V2m3RlmwkgXtsS4Px2/RW4QPbAPvj1ER6BpfWnPtuCX+/uNE0Sot1P2hYSqxSkrmw6+E
9tJdn1yEi4LKRAznXX3gvucPrzC90splMMqvo4y+hQQhoQhABM5u6fANABbfLCNSmcF4NTszeOqT
WWbmO6FqXmYB8l0GHLzA3SefRUd9SUh4gEZmxPla+rSMpIO4RdLDXmnwcWb7fkQwlfukQviNuyno
RI/qGlPJA5bxIsAhsdzn2HL0vHrhZfiR8mjF5ID2koUGSM2bZcqhg8o9NMm2npsBqDT9svzUsZM6
3jBATFK/WlV1cG3wrT1jIFhppOVgzlrWSDW5MqoLIneu4lCkQU4Zp/8dWr8rukc9cfX98OEe5Xto
Aljc4zV4dOrVxNkmIieSz9yvcirfU+vkq5h8JJCH+cjzJfPsAB1ixAKn5IXN89bZu87Y+2N0Q+mw
yZheNTobPY6oZ7vtOmcpzsIZWV8/ZSTIw8JJLuP9V6sJYZq52kU+1tMApCapdvsgQGwVBVQ+12x6
T5JyJvnAZHilzzkiLfZIGktYkBXSbVSGcq2rmTU49jxBSlQg7dtwCgc8NAnD8E0nbJrXDU4dJDae
h7YU+lS703bVHR98mqSSgc9z3uR0bKi653Kfv8m8pYnz65yN/rwmSIMQ8cPtJ9ura4XtmMJn7IEP
F8rPnq5DKJa8Sr70IlBb0c3QfzYP8V55qJtibqaAeAjaLAWXjoHU/cT8jgvBmFRO6f8dNDTGu6SS
3hOExPcEmLiZ/8TUX/Ko+4+9EFEiK0Pe81KUt3yHtfZDeyOc1A6tDwCNj+Nfi4FpNeuytv0fyatV
3dOn+LcXfzeUjDZMwsWX2ZMiDJBzLPBVAznbaZfntOmD/3TCTGcnMZYp0ytj/LumdpnA0SwlqhiP
YWko5Tm30nSIg2mkEwRVPG4uToV9t7olUjGpZ9lyskvdMtpr3yzqGv1+DiIYpha6vg+QWwLKMhap
9ASbsZjxT6LJlIGsfw/2OITAlzZ6exfESG1wLARJDpLWDwMTwWxdWM5qg35VkZyG29fyIq2AHECv
zI+N7D4qAl2oCYHoeny+YQr+GDuVN7wCBkei8XQG96PpjjJH7p26mHXBgeI6/PbNaa5Q2VC+CM3c
G6SFB7bJO/7iIr4bNyIqWgFRa/OfMBY4xrrm3saXkP+uR9fFuYEahyGWK5eUl7s5KPHnHbIbq8c+
xSHeZt+QguzDYTs0Wm6o/cLAi0NPm2ZJysRWBJUW3/2qRLO8M+lRnWN1vwzsn9mayV4yRFWRMnyS
VeO13YLMlohEDJGeEQlNxDO99E4DBIynOViqJc7hBhn9DUZiiuzrJb6avbj175104VDVLOh5M6dP
T67FzYW15RzV02xco8ydbW11qQyxRA6KUPdVWQkMPhtwUmSjhVo4uqQfwFsUOBUUNKQOYtPL1j8Y
qtMrM6xJQ+8jRT6TiUyARm2gSkgN+24n/OpAge9w2U+LHDtJbq3bXYCMOYd9zvj0DuHBmZXdLjcI
6cXu5q9K0M8g6haGOdTs5R10DrGs+jcvV59zIlEKfYiyWe9cTEANstQTnbQrAp+myacCZ9emk0Im
xA92ES+1ej0WexCtB6Ji7FRGkWartX+BKl5WPzbeRsMHdian6k8+Y9CT2eWRVfRF8uy7pcUMdrNL
hwAggryqAf7yaM9aiuNrzFGk6nECQwJR4hH0+OfI9+sWEN1CwKdS2l7CZ3aoxmD/Y0r4YccIGf11
oSmDXEJgSRLgCf62PTfYiCUmTxsH7CUGQDhkFTRpVEPV2l69hNZMMoCF/bAmMuk8CMYKzNVsNLDV
HtvABjuDlKeT+pJL5tVlmPFphwWZbxqgCjuePEL5mUgmJD98+5Z507obblIs6OI0jp8UUtuQd8XK
OnmKk0kcp5YYGDCRFQPIyND5rinjT3l7hBNpQEtimoizRq7DdkMEgkxfy8nIyISzuNqe/XlWAIPE
hMCBGUOzpiRRqGlHjUDUvIpWqAUB+cJMR6wNpwDPpiCSYmvdJI9KV8fhRQoDHej4jwOOB+YyimYj
1qBNwtIk2EGnza7ihRE1OYQ2tpjMiafMu/4LoTY0YfbVWjOhCEFItPqveBO7m8a9SkhNSjiQJ/bm
z01nwU7IbzrezoQ7/h1hQxxv9xdWQdQrhDx3aj+sQXQ1DMU5uxW1tM0m2k7ScCBirkWK+O3tTRdC
uG1i9/7pIsF6dWibpFVShNzsDV8TUkaf8FdRKBjXYSVyo5un6jYtCfPaF74/5k5pP7Crq747PUfB
ytwsSBXi762DUTluCF8ArCMaV/dIouv21SemViJUBHD5dVbCZcWMo+h7PKvW2vlbBUyhrvVbIQBE
u4cjsfAWYQaSfuOUO9doSyyKmmBAEZIDAIYg4SQF79XseLno1P6bSgOLZWkZ4YxSw4AljlvGrFpN
fsG5v5vqOMhL7TOSQ+uCrDXs0p0M7KkF9fusWcA9+ozPVKUKxeotgnc3qc/6lSIk0pZBWncoac0d
/Jkpg7M9i1gUt3nTLJbtCpnRGDzRFhd2wqxTfU+TDks7FBUcbPy3Q9epSJ2Eof5slAZLjEjsSMa+
rb7BDbd+YV35637MfhiMUgy1t83ucZWf6ZKRe20pJRT0O6mL3+qfRhRiVDAjFoL8aNmVtKOHY8TL
x+D210IB9f2qmvhtK2OqJRV1+98XHDsQn9WX9xbW9rWBaJro+He5oGvhppd+eOnxPTM2VWWMdYuK
fJNqDnFDZu0vUo4LrpIj1r2T81Q8ZcE+Wep1RIJ0k53J8IXgRytvGb4aWJHYyNYw33k3rmufIxAs
J7tsKS40+7WR3vx6+P7jAPVdK1BgfQRo6rN4GLAdG1uUlVN9VDmLarGk/uvz9PrWhKHLm3nF3aTy
MO0DqLrYRq8eMZRoyrXMrYqivvHnkSOYvik+1BZ73oGXHxOqsCBHq5oKyYjbKZOM0fJyB+WbveQs
uaZSdmT5r/5nvCmQVg+0VwYQ7pJw9bOlxNdZb4pbsEqsKAx9G40XdbeMJfggjH8tf9SB9IrrHIlA
ItSe9xKYEe2WARB+Z3Eq4/OGuVKtcXKsczAVKXkOYo1urmSlD3eSu7kMCMhRvStVa8lR+2jeWQ2i
yViW4R3iql5m7sOe4IBOkcirhpPNnXgHdNJ8f2JQ4Sg8MW/a4V5ok4I/sQBH52RBXZnr+LvLsiPY
LY6afRKalWNdlZFkwPUm9gHjltSw1VLomwYCBO5NZ6uBZt+3Wu7eIK24TfnqeeAq5St9OPtWfLSZ
1nIyfezqOPbeEwxXX4DdsgunhorXuXGh/W5L9t1mA27C/bxX9sQzgFcB+xM/28qknOG58oM/VfLx
V+uuOfWKx3GXmFhMUrxpakBMExEcgHA7QxbgmOQ+hcB64necXt7l4VmZ//cp55/5rjC8ic8DGyvA
0MFzl5IeNqgTK1OqeadXJewivHJ40GzGfs4ZmWfgV71H4WVgdjgPrZZSj65XdRDr51XxS90sMso7
Sf1iTbTpCsj3HvLSWIKjlvWPZla5WbcMaiSaWW97syt/JiPrI5CSn3UDO8x25a54F0FdP0GYdHUz
cv+PdMn4YaI1TF260Eed0xakqXmteN5JHtC9RE8qKEZ6krmfAYcwcvLupNjYvlnTJtngnuCs/+TU
eS/H8rsui0qj8QF09BlcjNjL70tdw+2mZJxBZGbmveX34p9EXsFpdcDyHijpfts7QUt0tfO7WJoX
Q6lS3goJt1ycvXSbw5LXLBHfrqEfuTOZEDeLqBgv/ETHjEyl1t0gRAGSRdnR8gscuJ91jAEBDhJ1
GUYXeTcrLINoYxJJNEaIugo07vmNdQVTP1ur0f6ZCD9BgJW/v3OaPCBVK765We85PWT7ZSz8EdHL
5QC2bMCp9g/qJxbQ5K8IzwlnN0Teg0u6SOGRqNa8GcAHQ9ioTt1D0LcwkY8dYzIThKS3lb6HE9Cu
Fxa213fIpFvX8DYc9RdToTa730nXbt6nrOeJEOdmuei1IeBlvRUoRTMmrOnX9U0tqcIrYoMlW10P
8R8WbaHD54vIpQhSyFs1+7uwqgP0vh+4oGgMKCO0mdXbNexfW7jf59J0H1UUc60yJa+E7eOC9LfR
TrUooFjfhBLBTy6Jx/ZLRk3BxqRaTHoGwIan5olX8lfpF7LZ5oJD9JChhhBFp7dCE3PQ0AmW5iqK
2xucMbS9af6GXCQmbkiuuaNz8GsGk/OgQwskfzm7u/th5tumMH8SSSuJUdA51wdFt1zX2GaXGePr
kLxXV/hobDMKlJ6z45AKZL4v2qRRtQc93p/ba7DHX3tk9SMZ5Tclc9fFgqErQlXT0NTlY82o//xs
CsQhYYQSMbB7hxgdkLKmmBwufs/85Bgy2JewwwVLIoqL6mLgPhX9J9tHHahkF7mozYUFD7U4jZ9H
FYdEQiYpCqczrgKEkJT7cNwRl6uZaI6JFbAs46XaohcAVST5F2uoeMkcvbvLgF5uT6Cn8AhC2WP7
tYeZYRnlUtqBJU6ivQ95cyndKGSsKbtQoUDyI5flDm486VH66vk25Xl+hwgUxiUi8Hi72LG59oBz
K7+VzC/cvvrxpQ8KCx40CrTriiQupN0AlJxlkk0xGeZsbGmon4UNkdVLctOAfXHX0W5cDGcsv269
OHYYudY1mBWNbsKWrW2e4PZI3hIU+ja5eFLGvdOuoR/ddzsxQLzXBXNgzTMxos0MOs9IekLF2/lG
YU1EDfuTt/UNmhJ0V7LF2xYPHJrCipeB0qi1MJTQa/fWvDEn/ExOXWeCtNNDmsfajGRFZ06AARWM
8ldkmPIygA257gtWUIcRp1Eio+wDg8w4fzxFJnC5u5AEU4PT7gDsh6Fdk9ZKm5ba8vsW2+Ildy85
6XrCB8OChXlyyuiTuk/yRxzufRv3hAqm4FNwlm3DYFTcWyrR0RV0WKkJEzMUHB82C6n3CB24hyuO
KGDU+G5plfTBVegKulEIlKjU8g0ns9iS8lrDxuaEgABlatwqbUT9zavIn21kzHhzcZ7UZmrhrD2Q
5FdYWGALLQokdM88Fgf90CjAdBLHZAmBXPl8glke5+HvNky/7X+w9+sJoBlmC0QdtBSPPOGx2hm2
PMccbeiQEKVJkYjTkECOAUbgF2Uq6hYBGp7yhWUIJKjKrzrW9hYcEmEdQFm/H+BWF8FGrsEPtwJc
6xdapsWSDYcbxPgt0NQ2FoFV6KH1t+/G0zxprwNCHdzlH6wi4qJFwROvRSJhEocrLNmHMyLue/fs
RbnPmqPt990uoYU9RxQ9vwyU3jsWzu+897slzmJYUXugbdItzL4W1RwJypazAy6C2srpW/lfLZR1
Tgu9Y+00YKqxNEQd7iynRLc+KIexwaF/ZJA5wkCJ0ToJ5UlPRqeJfqIQ8HfDKglVjZI7kS6je9lq
ppaTUxunFxTkqWsaJTJHnxakQJkxNm+P34XPFzgcOaedmIZSE1nRxEcEx078GK8sK/byrrkLajzt
EvISJT8jWLNrz14n7MGFE6H/TCt6nKMEewaiuNz5P5Ucm3ma6DpSfQKXFyiJeX+nchJqDmP33cOo
a71Ibioz2iOCfjiHEUwelkjILUmtBJ4Xy29HPCR+mKNIpPa+ityGfPxlJOvw4gT9lNzawru+It9E
gRhnbNpoJq7HlYPAsj5wfKL2WCZDKhjJGNsMiuKLkpewGK7vNGmX0pA83L+jJWV/W7V80Qci4jfa
WbTGE1rIP6bJd+BufefyLHPKz7swdIZoShBtPlvDZzm+wvT5hpQauV/F3EeulPKgO60AJrUUp5Gh
U8Ewa8YdO0ms6GsSeAu2dKdCSc16EtlKP+HbVZjVL88N81cxKPmrufTXlqIU+Fl6yRlAfLRxvubQ
cWjzoeAqZFvIUXvNZ+ujRhuTXkXgDy7VpUYThY7csfNQcrgp0KMSnfJGApTGYHUrpwwjCdiKrWds
7n727V7vKtVRBHoVLEzItX90yKnjC8TyePCYQtSCYd5qRcq9x6Tbj95emm5EgvMeXSdWe4c+twjN
4Gyr1j7nblPGF3ZWWL/MyJU/dJakzupZRCYZd/jxJPo/OyQL2i60oljyx6P3ohOGhwhJGTpce2e1
lEdm6t4Dl74uCDqz8E/jNBk/D2tBzs3Oz9Jshh1Js5w0+J4HYFoiDrO4rvtFJCLt3fPJlyDhua8v
7oYaNxvetq25QxSV0lQtVsQCXaKK0cKAEB6LdMfp0rmJGb8UQ2PG33geK2IFRr1uif+44+n8ch3o
fQbSJYXUAJoL0pYIITkG+cfM3r6PL6v6JTcbUu7cbqvsPdx8UDzu3kprj8BqIoAEAzvzjIhXl1c+
2Xjwf4J/F/SHcF7BDKC4CAlZ8C2ELs7lodrQtoLc0BohLt0FuVfBvUjYzWOQ7N365/sX3DNeG/gz
1ME1eUDmZXJ5h0kEH/PgQC96unM=
`pragma protect end_protected
