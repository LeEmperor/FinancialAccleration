// Bohdan Purtell
// University of Florida
// Description: 

