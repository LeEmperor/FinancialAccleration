��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��x���9eS� ]�_g�Xh3��1��63�A�1{Վ�eb��9��d8_��g�G�oWs$㩕�䫀�*Q���7е?-�@�Z��.޷�0�Ȭ�*
XL�1���-ec��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��D��ÊC]o3>��FyM��쟪)�����_7�Hޜ=���㗛�s���+/�d ���e��`�i�'Z8�gU��̓����;�h�9r�Ó����sQ�35�TX��=}�>�O%u�Jg��x�������;S����wI�����y��2 #e�d���*�Q��
!X���}f���S�Z̏�_�d	�c0���;k�@Q2L+��ƨp��盶�z:=JuQ�U*h�0)�t)e �0�xg0�,6Ŗ+1>����]�)�])�t�ɲ�#
w���8
��$v{�?�=ëλU�ȴv���/U�V��Q��"���(�2M#n��&��H9:j|w+k��3;B9 Ѣ��׵�#ɡ��T���-|Yøw����F&�j"Q=̵�\.����tnK�I�9�W�9�9
h�+

���+F�2�1
�}j�T�b+����#�ɖ&7J�nhd�=�N�q�L�u�5�7���H�0%s�f����W�"�e#���>i<MsPH�V������6�>�)W��������bre��g�&�rvQ��+�(p��c�
�*G53��PJ����ޟ�my�<y� �5�zt�j�m���d�5i�g`��n$�9�
M�C,�m-}lEh�[�գ�Y���mv�8�I���	t�O�n"�
>��g����{w`�$Ѯ���5�����h�\��ay�;���_���Qע���'n�q�'��S��Q�E�6�h�C�M��x�>�$�U4Un��F� ��//)�2�������1�w�N��*\#�W�B�畚!���V�c����z)'�4_���(�����*���J�St<��=Z�8��~�Jl�r�wׂ>
����'��u)��Z���j��Ք_$�&��'R��8�����8%JFu!���Vt�@&�\��h���qQ�Ğ	�vNbi�N�*���b&c ?��uPK��d�.6�'�D��[Ho��Ys�-�x���F�ňs�e���zmPK�i�m=���}H3zo-��_��g\щ�@wk`d��[wP���^h��HۯrH��r�稒�uS���M��3o�� Ha��������[����0n+�;�`;�z��>+?[�� ������h��>�M�@��p�s�h�
u���~���I﵂�YPLW��;1Q\�f�\t�g\�\,��l�`��?�S����B�I����~�*r�g�,粰|4��Vq�s��F�,�@��� ���ߧ��(nv������b`4*v�!>OYy��S�^:�4&s�=���R��X���?M���0ХT��Q��_�1	/�D?�	O���ɳ�N����Oi��>S).�+ޚ�8�n2`����u���Q����6�3��lNՔq;�r�J͛b�V%xp����?�IgCU�aHϗwk�Z����
��̷q\�����S��*�ʶwHk��7*j���4���@h6�k�����8��c�1�q�ɫsjz{�/tΚb������/��0wǾ�Sw�)�~��ͨ���2����!^d�,��\���H6`������¦��.�=�Onn��p�G*{���N�t?$�C/b/�~�MBe��xڀ�H�1x$�)�i��o#D�ƚ�T�;�Z�=�p��t���o� ?�@��D�}�_0a�3�'͖��FQ'�	V���P@u�r���?H��-��p~��F�el�tAvi
�w0��y�7a��)C_[�fa�����H��:x���ZDu��y��jFjT�	��q� ���2|�FH�l��� �K.��6��2�n������2�'I,*����o���;	0�ًx�]{�J�Ѩ~4�v/*o��e�l�v�!R"�9�g^��h�̱�����	vM�p���d�u�ډw�5o�C���� �i�p�iU�s�XV���! n��5��ΈA�YCCr��n)z�&�Ln��굙䊌W��^��┊J%G�����h����C�ޘ������:] Ę���^���ɈUM�̼�5pF�h���5$����CB����e�>�(g"�T���mܱq\��(�d5����B3�]hs'E����m����sݫ����\y�ݵz��V8��X$(9�!DR�L�1Q+�%�ig���[�|
$m�$&ڱ
�y���uc��h�1�p���rT��?����+}�G��Txμ�_F�ȾE5l�C�ϰ�ʀ�;T`OS���	)'�
�����J�L�(��Q��\J'��]ƃwwG�.�ֳ	�:�0��D�J��<Y��N�?}ޟ�E��K��������j��(6��{��q�p�Oپ�HR�gZW{���6��т�0������ㄵ֊J.Rn
ב]��}pG^y�$h@���� �B��4"�@�q~�����;�;�N�Jc�i�Y�vRf�M���J��]��W�����?H㽠����9/-�{�V%�.M��p�MP��p?#�k���j؆���CL�BK�����qK����!3�K�z3#�Eڝ�.CLc���{�̊�'2wZ~@��O(������UDې:pf7mi�p�K� V����>��w]��R���/5��='��_�'g��j;z�<�Fm���)�}ҩ��j) �cՖe~� �n�����Zm^t�Ըk�
�.����T�g������UL�z�ap
7��dHV�ѐSN�* �q} 1�<�#v�2��2wM��~>�U޵�z�i����,Н�dy�9���(����p��G�XI3B6]���3f��j��4��م�,%�,T�rx��#��3�oϛ�C�nү���_�|�3���
�i��y 2�1W�??���I��Y���'7v]���={;��Qgg����&c���u�CĪ �f���^B!So~�HS1���C��v�$�>���V�C�IQ�
�{94��Iͧ��#P��h�R��LiH����"ឃ��f��/Ƥ�se6�)T�8��ۓ��O気��%4��6�;׊��So\��[j��T��j��X���'g]ރ�X��{�4��u�Nđ�fZk��W)��'_���� �y�e9|`m@J�|憀��6��t'��#�L�� ����D���A���6�|f?�~�QD�I�+]����(�1���N���n(2|��}q�dGn�*�YC2�t������)YJk⮀���Ul����۪���BC%Zڂ��\��*�9t"����0���K���LX��?H5Eu�+5u��� ^��e_�n}e�e&׾�%��Xl;=�c!(���{I�^ݺ��^x��q�������|�t:1a�؟�����_/�E�d�},1�K'8��Dk��ϼ��x�{��~�Y��xч,u�aJ�<���Ǚ*��0n��$@�B����1n��	�f
�ؓ���T�����#%��Bh= نB'H�I#�G����=ѴJ�͖����'��^���>���9iny��U�����Z}�� X��)��P���]�<(�^�
��kށT#��e2o���YJ%�<�R�wf�-V�ʴ#սo�+��I��k4��i�l_'>����M�ޯ�{�P�;�ݵց�fS�� Y�Hbڳ�[M�I����G����=l��Ĵ�bC���l@U�������S2(���O0��f�7q�ٳ��"���+r~'��0��rX��E-�բ�3��+��ԝZ$�)#M�0}��A���qī���ʌ@����:��7�0�K�e:S��\�t��j%$�^؇[H=�~8A?�+�+���F�� ��kr��	3֦��17�E(�"�V�M1��u�����C�rE�I�b��g(>�5�� -��#�,��wo�j��n�����Q��Bn��HHayUF{�ݬ����J�ߋ^�\=hT��ޗ`�ɇ�j6V%tZ�|���N�3�4\R���+J1��ނ�����U5�W~��wK��k�N퐖*ڿ\�.f>ҫ�>xEE�ݓo��Kz�,y�xp|DD�N�ˣ��)���vϲrb��,�N_*`�v�䶴R�D7ZsK/s�-p��ݓ�䲥N*�!:�?ɘ�#`1�,3|ҲŖ3qdw��S2q� �lQ��d���\�IsJ9��/I�������ÇP��3B���#�����J�i�71-~���/:g��rZ&��zQp�&?I��mAr��raWl`��ڨltͩ�ܹ�s�x\9m���8!
��Բr���Ң�V�i�$8�^U0�