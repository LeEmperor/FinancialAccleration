// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 19.1std
// ALTERA_TIMESTAMP:Mon Sep 23 04:09:48 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pQgQ98sgqVLgY/QJe+KEvEoU1Awe9ek3pQ7d7OXVa+9YUbY5rXC4Odf2z6EIzwEp
vQURcJ0ThvY59Ku5JNmL2Ev7U+/D0KO1UoL5Fxx1Sbk9wnJNzNhOUZ1tdquj1+37
2tSI8tSz+TGVK+r5d2Tb3bUYAhlPtac18tQEp8PdoWU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
+4AJZajpa9OUhIabIYU5QOTBpdbxVIaKBu8czFH0C2cJjuAOPiHsfGhxsbr7Uihs
tQeyn6gQhiANnZoQ4FA16ausQ6OXi/2HlpHTqNdGBuBI/PBQVAMCvnYyAfJAYtfD
5gbSNV5Z8D5phqZM+jSQmprJfncDMcAG7FCsjHB1OWQebGbcpWE0sxRqEAglMuKP
DdKF4M3L8hL4eU0XP0x5fYGkJcwPOxq3TDCuyuqk1ylMkzXQYAysht1JQ8U26oEU
PZ+PEkgsweBxcmi8fOmr4L/4CK5Dap9bD2nqlj+b+vBWeqKK9qJOohvA8xjxMQG+
w1IIPnIQDV6mpyvZtDg8sf2u56f56ApzTs2xbI4Wi+0YofXegKu6+4jLghtm8S3H
6jVNeHjFqXfB6Se3BTHwCFcYs4WkU1C9tJ+zo+S/a6wSkvvkeFfnzWSxGuy/BnH2
1HKEMTKKl08HvRB6RDM4Y7T/yEYfnURUNUPHwSW8zIxJgfKpnkrFrrLf1a8IN27R
a1T2o2TgISQ39jeYEqJJyJhQ0JhtMb+RBGoK/Ouz4xSaR0M3qve8WARbfBlhPT2Q
9k8u2EXpTvwDjqORibpzHtCTRbC3j1+Nm0O2QCucQrjUhpDUQkQTvdGkVcErRRKs
n6clACBxrc5fjDMXr/K0AwvX1VkAgYcs+ELrAF7kH+uVrB4FhV4uOjQSduIVi3IK
2IOfndd+bmaXUaifFlVLJxQaFcvHa8B11pfAhgn4htQ7/I6sqWqu6neOXJe55r8T
Fyq5NfMSMjLsJkeIaPiLKndp7uKOJ+w6vmocbksGYJbeWN8yWSD0EJIlrfh/XANE
z1fmr+di/BR8GJwFXfmpAOeA0fMubSeGMpOFKH+hF0nERNV7JNdnRLtJWY5Q/d0C
hMuV/Cwa5EhfwFFhNlHGe8uoxprqDM+EMIFr6EziwTyiPg3UH4Lfje2/3xAX3rVM
inhSle7oQ/40AhEgetZWVEkC+Z4jUfq4vItyVvUN+zhEwI9no4qBlh2OtmoWiDVX
3QV/uj1qqPinP8Sarrf6J6Axl+es0SVQGZQduig3jc6nVXQ1FQqd2TdhNAZW+vWa
OGCOVzBnc1U594EGsnzL5W0x/aM/75Y73OorqydHfM4yjNUkN+7bq9hNY3dCRSMw
5fL2ChNCi2g3d0324qeP44JXwy+h8tTKv65FN2mJF7EVj+ygtL1vvA8VTe+CzHoQ
UUBvqXkLN5Hyw+mG8Si0F0Wkm8OSq0uajIbYfGw8SN1BH86mtCbZcRixFFg8PN0J
sTZZM4xLQ5lOMq2k+pvKw9euX4HdZlbMdvYy9x4eisowFBFbZFaG7ihKcUPuTSUa
WkmgIAPXhY5VWuSZ4EhVK5kkvx5dzNmd3wfdhdeymazqFwC5bWrHIlwMztZ+gJRt
lPsfuP6xUbsBzV+1OpllJTeqCg7IkC7Ea3oY4R6iwN/Tdskh05CIDcZV6qu4o9zb
8w5SzZ1hTxoKgSRLBCVvVTuau+5CLcdAv/i8vJcfG/y0fd2MVcQAgWShMoGE64T5
ipO4TVCtFygI0M0UFC9E9qv45qiSTRsww4LyxKVJuEB/Tr5AbKHynlwomOQdffon
LfdyNE1g1nPDem3v51scIjRaO+xGleLPNNJi/4+6f1X7RGD7BrwJySVz1tJ65Zi1
E9EVvFSWyhkXTy45FwYCfuu6arRoD2/VSdZEx+md+qs0SPN6j1+F8xwriW6NCnoH
PqG93X1eDcj5XIOm93dldmgzIs/cCaNmFSz4VRUaG7hg/OxcMK9Hzhb06lqIq66D
ZUZbIb977SMnuONcrv/cTUOXbBW2GegaNal/cPwsF9+VeArcZ115JIg5B9QuE/Mo
AE2ynGMYbwBMPuNpu2OtzM9Nd0UmrgkSUmI4qHkf6o5Ii23AYdsQQ4JKdze9S4R7
sjTfLCAusk+btsCAwuVi7vBE/rBdzex8zsB7KrVyT8dxH79UaBm0nlAfgeKQYRLk
tdRzXP3YWUJZRyAP5Ss6e9GXdiTAZYWpAe41tf//vQ+hDS3qjH4VpXANgz4y/8+c
OYjZC96QRraoOfeXYBVBz0hCMSVnm+nWp1w1+YEA8qkbMc2F7QID/F3DpFFSHD7X
BPLdFDPFOH20ljdw9MmSNPze014WId/y0Ja0tOEWDUph/ma8Dcj0BqnVmgRto0Pf
4vNRwKSF0Cgqv+3MMPP1iWk4jKyHOpwzXTKxo1SIvtjDdOLWJ+HPxMGf30R3+jo3
jkDTp/NCeI3E2Unvgfwxcn6HPa5a/07xoGVuVwMrZo3PItocdnv8Q+z5DoNKHy7T
FzvgkhtfyHYZ+h6piLBtHvW9F80zSamWYVk3+UlUoLO+Z65Tsa17NxnKnBk5eePq
hh9+vk9pTViyDDqzGcZFv+hemzuIGFOHAK1LiUz/ujjyclfzaBonmS6EMnpNByVL
ic1FCZ14/K2NR0zSDIis3FWPg/zt4APucL0CIxJFpMii3BWlpRdSPl3bk/wfte4x
O4u1gFr1CcrJCZqX31Qqfa78vG0V+hA+JrRpvszFvfifaS+yMCrPcg7n78aKxSyn
tl3d2Kt9UpSRjewY5UDGYZkGWIfokviqKp3suxuseJWa8yeQD5kP+0HkQ3YODAAt
y7AMrlZ3hw9CG3I1O8MeWRevwFzqyWiRc9vDDy8SNxx+3mmGOj9Mf/KZcAsDg3O9
BxXk7nVF9gfTHheJSDm3dvThji3uOthMm9ceWg/bwAwNDEC/b60hwFJ6WdQs2tOj
K64UIfcJj22sBkZrcEnQZKiYsxoCPPSMIgGX57GW2z7htbU1xyTHvB9nJsegNaGb
1762Jzeqts9iOMOpvC3I+cltZ7RGHqmWBk0RgkcCJXArqCEeFfsFhH5013TxvwWF
kbOsWH2on/p3zs4szNt48QIUKylbECa/4cTq2EWvn1oxfZH2pF0vWpNG1X2b6PYO
vslK1PH+Y5XTKVPfW1ib4bn55Z7SqicUdSG1TmwLFm5eHmYGWRDmg+nD3qfCtJ8g
CIEBJFzfqKkFudSF8T6g1C1E8qWQmMtp9BnbmL+fUQJfwNO8OcU+LhRl81OLaptE
gPD24c5qOTn1BEvnJRayu5DVMUlP+AkwnYVDNQViO434p0bpQusJqu5aOSsitLug
ihHLty0OJJI/w0g8bb+NUmvPsKeQc+uE2/0sYFdqXmSStpt997Lce5UyhJBijiOS
0ORdWMx34mGG+GN32+VU/ks2uJwgM5jOm0KFgH1vQPtVlY8aZrss63cXwxy9sqAs
h34AtqIWRBVpEcvQ9pCEaHrL8L/2AtnkwuVTft83ETx/hlvi+haO3B1zB0WL8oVZ
M1HATXJ616RHjZUAkshWLU0lIcMhH6s5019RYwal0rgLmK+mlgl0oDIG135GaMtJ
hh36iKlEtAEhoEkYqZ7OPSweuPbcx3IUgi7J/t0PhX2RSJw8p7Dz5izBupZCo2lh
LyLBk5lCXiFZtVu1XwBMZn2xCHSMIYJl6RxTPsIrs+h6LZbxKlK1BcGWsSmnJGS7
hk1XDk5vGmo1JLXiDD4vS+ppowBiNGBzLoepKc5eLjCK9ChYg5d0eavAzWDNddOJ
gAzJN12m7rJognkpszBfHbZxLPfYdnCaxFZ8F3u6JHBWrP+wE/XpyTibGzGBa7SB
+XXM61fbvtmZDSWDV9SrbztrGGTqz8xWvuou/R/hH037irPj4xJGBoZvq4Kgr30d
NOW9CCAUm5HSeAuZoLWxX9uyWlLK+8WRHVXC1HQDmoMAKbQPqMF5UQJWwSH9INQr
XmLKtRJSeQW+Rh8MSt69y8fWlRs2sZnIGc27f1O8Ztj9g3QDch4XgpSox2G593E9
UalowQN9aEcJ2jR2PEAOkbUmSGv8Ewv4ByqfBN4nf6ddEhnn8WIcozzxLs1bsXCA
dNjCedUohHpcBmNex85qalgooj95LAvFXe8vPcWQz7xP/7ewp247kH9J7QAMTkVx
y3PPRbHX0SgoYGXN3+To4345SPQ0Th7R89aA/9REYQJr24BUqMNFkMisYmaFXTln
nNWFDjUSFDrFmdZascGESumtkOl66u3yhSY18IyHaBY1LONoFBzXjLjAxLDAV/Tt
l/mujvVhokgb7s0H2wKfAV/WNcepo5Jp2kBjckjcjK8pLU54q/fnFJDHIpl2fWy/
WvIoFq6EJBG3/cwzD6Wpb4/83phv3rHlLje+PQPHRO8eaRwou3IUJvjLHvIXcrk8
2A2rhY7tD9Nsi1VRpoom7nP2pm5YNnOVlmCnWovn1E94hdiTsEtWqt72Oblqcev9
2jDXNOcO4QOQ85cDJIf3xmYB8yscjsPNILb6p+fdf5snAedv72czkPdVfCRuRO5l
uoIOjza/TQbO0ZmXc5ZGW8ONB33dIPBaLG7VpjPGVtgPVaPeikIrs7JiXzXRId+9
r0WustFClHoA+8mpEFQxZ8fqh4tFb0HCq7SeEwkFkmrmEaW3cbWdgeoCqiNOUfPP
XIZFPe17ds0kKGUZA7DbDuYN62ebqJpxYe6zQXMrniCOji6arAdZ1epU/dzPejQi
OLM7SZcC+JDnihC0854Bq7RvIW/jip147VCx15wlyO4jrsqAp4nK+Y400AERZTfL
0ADHWpuSYfu2HYIA7M7LORifCA4gf+aT9HYeiKvRkB1DnSb6CZrR5aOIiD+bqdag
dk7c8zzW+G0vETQWMf6hxLCwk9Nk5yz+g/jeWecVS3dQL8pw11hoZG1osINLmWsQ
ncjE66cS323U/9D4hsRY2XVrv3jp3Sg1kriT1WkKvXUzT6G8MQzjTai9+o+XlHg5
yPJO5VzsctSpJv4wfHj9YDM5wZTgfBHmdN02NUhQNiyfLsEBWXrASFW74At0BDgE
DQbWTdtyr7GBwU28+FRBxK4yTAKiia1KjasZss67rgHr4IcqdyYTjwhBmpJxZmOw
Btm2Yno5wgEv61xcMBloFz7av5CBmqNsV96jFShfu4+0ZISr0d77IMfndueraQE+
U+0EPB/eR6CH7jukFu6TYKTeoa+Rq4mY30lhmpDGWuKxDK0DBdWQgRjji017jJG4
LJU5xAdxA+xsSRDwmmaBMjjYX1EdcOsg6UIqj2pOUQx1eKzs8RnkOxFmf22T4xmy
oebsSsuwvDUm2mXRLjcLdWDzlyeEY19SFsneiOoRhVpBYDInrj7hy0v2JOHpAk3D
b2O8zd4O/VGPX2h5YuDxBZ414ER4ZT0eJ5N0t0hrHAtMzjiOQPOZJ/VYpmkXPL3e
CfcRmRijUSujpjg7wkHS+YubJT69I2nJ8hbh2Y104io4Plo4TZtS/CkZYS3draUN
t5Kf4H0sNA49arXVQfbW1bXe02YDgNUcK9tiJu352lnIuGHKRKj+SrzDuAgRaThh
oSX0Wh1luyyqpnB4hySvDcOEnop4jso+zR8pR6J4K1WPkHPTdb1AikaPJeirshzg
14KPYDzgUkuLK746FUK//2/MrHAi9Akzp28ulXcIDpQDWiulaOVwOKUARSwypJ6R
rB87n8Voeo06qLKlokWkObPPDb26Zh34oFSITeQhXQy/DeiFGJS74zaWGv7aaYIO
5uf9d5F5+v9FZkTG0lCEtGrE56FOs1u24p0ANrWKP4jKpPuD4V2bPxp4ZA++aak0
32t6GN9akHrenQlkymyZirR9FSHDjhYb5jqaYyIWaTtQ6NjZegp6szwHrx9cHTMz
r1l+oCWH/hzXqQCSm+yY7IkvDClQ4FXdofuIX0hSTt2uQ4NY5wyCcxzQe9PFX7Ai
kwsPioGrolO3uIz8gYelUJ+v4A8rDdrHeR8+jSpFkANsWEVy7bXyu6tVpw0pJHiz
So0ytEtY/lucjcSYFRcvL/juOY5UnidnGTFlCVp38V9h8rOA9AYbP+LCZFVHt03U
ANhQD7A9KOlnyItKXakHT3EVrtWG2b7KjU4UovGtD7Mpy3uhS/kHMjlY7Fv48JCv
aENtMMgD+mnHcP35g3vdxBnbdp7XU9854rPnRjMCv2YW+vkhYE6EJmKcsDG+ZPMb
o/3eKyzFR7ODXFZcPJUS1t227NtHaLCBOmwFFsXZ0NQGcMKcQwTr6sOTkFer4CkO
gn2mABEvgZBTfcObpoz/ACawTzeE0/Ugevt6eRJn9t/ylTuTosOaJMdZSBd/3maE
thTCRvhsbUzszoDRlt9Cux0hs/fV3ZR+xLmmvdYVp1G8tm5i3zqCsdKDwPI7pz77
1La/8qAgYCHtGFP9PzPT2mfmWtO2+KePDUzgzSa/0s8nnhZsAlQY8IdfeLiJtobS
kOEtsc2w8vZNAyvUOxhZcvu98QUYJ4SMPAwMvNLuPFbLj5V41jFqN1fZQlxfTPEh
lVNTSbxW3Z1qYftqXYNq8IO7tU9tUa7ZC7PKOf/hkPZd+i/fsyUCw4uKfFd+wRE4
2njpQa03iHTGn8fEl6GstCKesVcvshWFHrE/Pmup1w8eH68Xmx78vyZ2kk64jFqJ
FOBg7jKPxssHOl7McjddtYMl0aLI/g4UctgoDq5KtgtG/xrvZ3qzBTDVa9+qNpQD
0e51+s5zTSpZBu4gU+d5nZRVeI7Ex/ZfbyUKUeKqJhF1GYTY7dcaTAlVobdzDB4b
imnhLC9IvMlklWHN54LVqXjrFeurOQaKLFyzdczvNmkgrCyJR6ks9k6I/3v9NU2b
2W35XM/YKpbs5LSSsBBw+B1bvIHMZCJvizEWMJq+Bhn/fgPj6ijQFT4k6N9sInjL
zFYRdh4gRoDSgNp4R8ghpJadIYT0vw8u3lRJ8hNpAdzBQ8FMpl+zdzx3mGwOfRsE
rXZz27+QlTBSS2Om4laWmGS5q1BfoRA/EtKxxBroy7laoGwquxvl6FBzcXqn6kar
oZylwVj8DBsfIMGt6wm54c3JFypKD2af/JKXUImObAUTgQd0aaqNKwXgT1PYKjfy
YewY42XHyV8PwMxHjvsnf99R6JMfpq8UvZlpAlkbjl+I78EZzOaxvpUU0eddScXb
FlOVCLykqTc02tn1F4Mcp4T1pqEErZlZ0rckbVh+8/P+z6YjG3f0l8X+F6x0/MMv
HzvBgDI4unEbCqPMulR495BSKoNzdv5ySty9UbemxXI6r4gm7ttdAhxTIOMfgWs2
WykmW8GSEblCE0UC7FThG5gL9TXVGp/Sdo/9/xZyMfFdGH+XSqFRqhJ5ZPagiBAl
1coCXW1wTZcjc8jK/67q6TqGjWEF6DyECHzmFLkGmtpxTmdOGPC0NQKX0ZZIrikQ
NY+T5KxZiR7WfmvtYJIBlFkkq/05ZMhxltzIJ7Ijd3+xQWB/HaBG8xkQwSic+VnS
nkiUms05oKILuQFLghK5HVWIyhdncSEvMziIFHWHv+HNvn3gpm/CtnuXaTkhSnG/
QxJDj+0In2cFoBF7/cPKTgtluwJ3fjvj9whIYPhwLEz1nyPdzLFJbLxEetpILxh5
Wz3nQp84k6n8XTRe1PhbJnn2E8wJGcOdUly4A3fKamNeWm5mNZP7emoVUjr/EA/o
2XVjrpoSU3quqBEuZFezj55lbjVzZigEV+yrXEE8xGPizf/6XJtn3c/vM/NZnUU/
pSD5tl6DYheuL37O26hyyhAILB3g1RvRRuuWRXgNa9GuUlQRgKUX+eLDz5L67KWl
+1O5A8p89WSx+IftUICYhTRlJvnF7SfRq3QSRe5zVW0uStdMZ1/D/PGhkX38aaW1
5FVhJAaFpKtAcJ+g58FlkNctFbbl2R2+8iyqKgc5q8NUasVyTTcspscB6wFY+ErR
re2etf++zyluYsRHwtw2PGd/B6/YNeZlGqU1Z4KgHKo=
`pragma protect end_protected
