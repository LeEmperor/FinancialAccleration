module toplevel_v1 (
  input logic clk, rst
);



endmodule;

