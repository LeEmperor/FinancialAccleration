`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HiPoSU1LCyzeIQyNy3LHQY22dIV/87XEOqWRdEJZ7Omw04E2/cnYsyx0Ok+/hN7b
Mx4Z1VtnFZKzRk1LJ1UwX8k9rLfAkWLL0tEV854QF5TP8ZtQLp6r1Iz8KNkw7UPM
pI30E/VIlTBZzaNcMTcFpBaODrx/Mk1cknlIYa3Trbc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
EMihWJ1g3V5CAGgd8HwBd0wlC48prF3a+GQKQNj53pFsN45zAVDOKn9u9cyQ6ufg
qI2r4vA+OPzIH0MndGwyzeDH9rwVC2SA9dxQ37kN3J37rM5wEYSTzHHiPSNMWJiQ
jz5Beu5aDUiYF9Yqyk9c4Hpelsz7b20+OCRNjjqV7zlzSVLwnXw5Rszt6M665y7N
YkoNFsxKkykePhR6PaCnG4vhEnyhpPJ7t6ilTnD6au0v8HtgUVnvX6BVyM4ot/Eq
17udTiMwhMRplpqc3Ht5TaQwpWyg2dPwfqrlxtwqOQyFqVTCfj8mylndhdY/uatd
LqILm5WDkMFHpH0q/q+twL9mJbj0igtE75v+bOO5oz7K0Ob5kqH/CaQ32+vAvRhv
4Oc+BfJ70Vqq1NtI4ytRMmQcbF4XxwDI3BTBb0LBMveA1/jB1SPSliJ6PMeJrhmZ
pz1U0gHlJPx4Fr2P+ziUFtOYvMRmeE6tr+pqkp1JOUKWUgtMXSo+upm1AhbJAs+u
ZiidyJrCXL/c4cOQ9oRlj1uUe8U+juJXXHrurrhSAfEocV8Ageqj4WVbSR7F09Gb
vldaTb8IE0CzuoECjAh+y9gqE2taqbWor4r3CLfkbw/3I7LZMXv4lFNcZ/TTzii2
ADhJBJqIsHIvPA1QSpruHm9zcdZ71Xdu8ZS+M+EZAt9CXWFYiIknKmaM2xls2Ub8
kqFZR6+5hcUS3YIBRRll9w8S9MqaWz/ISz6+018ireaCfhN6Lcp607vUyivDrb67
Xi07s8QHRZVQBIGzRG59a8/X3od6+Y9IQ9ywL3+oBTdOwl8RszBRoPteuc42qMpf
1QqehGZfS6RIfw5aub6F4p2RIsjW8AFnZm8UzlTGit47PA4rwJU68LXNB7GWh8uz
pREc5oODFWz239vcT4M79kouLzxevQiWIqSAF/5woLW10plSMH5Z+P85aIJ/EPc8
OCPxiJKcLrGSp/eSCDicnEe5A+tZo24pV0XOpgg831UFSqUBXET0vaUptslUP3ue
nXwqOFoBSUVn70PBkZbTVtQciaEjoKqdqKyHcQirdAii1IJNQh8krnvRB65cSn4X
rwrp+hG0IoNUC1bST8lzSlcXjX8bhxDw0z5NMLp2MeEuomUzmJaxretZTHAIO/Ia
FkJbFky2771HETCZQ+l4IC0rk24K2dpuTaPWtJVuk1KsBzjakIVmaKXZJPAMeg43
LIbrmMn98RQFbyrUau4hcjXdStZhvlV5hrIzz0P3c0HULXa/PKEnHKyMxDMmDItK
Patgokrlx3T6shI/C29/gv+JYpdH49GqeY7Hl076RwQYehkrRwRGzuY/SJbSVmH+
DMh+wcLC/Drm1MkyincrlHrAqlzHBBZTzc/+tl3KGodzGpUmV6gHtaYE01MQBy9k
hIsvF+A9G0cTB/mDCFxdD74c9/7nlCgQl+6JSKXw1RUwkOrCQ5zYsHzHz/8doNdr
9hqLNv/xhue+brlcmMMXcO/4KHABh3Uw1fSPU0Y2ocr5eUFnQtPZ1MF4H28wRbev
3R4x/MoYJrxA4i9+Xfi5309lKC9qRIxUaVlDZJItN2XLwiipFxnPTBLTSNs1eozX
k5t7o+gqxlFTGveGzANlBR3ZEtErvpfWlFXpBcCXEeNelt/N8ozzq//QcR235MYj
1gKR3sZ7otlXK10ll/ylJBdOoP+iIBvCwOfb7CeOHPvzS01lFRx1z+XwFsGL6LH0
fO2MMeIMkL/DlzjrffXT8id8JhUfsi32U1YeP/eIlXqWwCnh71wNmaS909J9c4Er
QBDsoX5SE4PrAqvzyCaYqS6m9RVUWNa1iF88LbNgnrpipbgyi2K9xXgx9akoOBfe
3e+SuFNRe1SFV93Nw1Qojf0AtRrfzTKEF7UwK2HVqNAFgg5eK+Om8SI4HSH37S8e
/DhgfJYo47xLEbSZaqAJWkdtrpoYqkjDkk/XEExnILiwyJZKzQD1QMfzYRSSylRN
bdTOWSvFl7DFKN6FN0FI6XntW/ZE9Y8HQ9tVeiDKxdyn5q7S//TWSOJuIi5DFOUN
fFOI7yQG4QNexQ/EwSlmbGWJ/Zoon0cs4/4w86OR2TZ40dLi0RBivi47IpM/WlSy
DdTe8zGBarXcamkKqdpRcMUAzNrkIXD+3ftMhGN8nQvDfQVuHbXOr0na9KLKQqZK
lTyJJ4GQZiO/1Wsn9mzPVGBOyxpIyoe1udypvXS8ptW5IXUJ9VSugrmCMw5VuMk2
LMzS/R9UjfnA+tHMYqE99s39lMSF5fBsmUAPZRvelW6tOfD28CIBkZo71ADQgJKV
exAwaG3H3e0eVgVfda0E8cxOKxw9XYcjBbMWvQOhL/Dwfo5mVQWC67AiFAJm3npy
QI9SJKJm71vdgVEx5N50wDSIbtRNWeur/C0qEBVmjxWLpBIiURx7grToyIaAuJA8
qBrI88OnYAbHscG+a5GoJXiI8FSDzANjBgzy7s5ZdVFGO/e9yfsjrhBlIhxYsnO/
AXQu/xa7q9hDWkYyF2+uXHUTMKhRNmD5/+KaM7gn6+dEceog5RW6gL++lTah/Fw2
wGbrPErmSGhhpmuoPRPIhvuHbeiP20pgqhjQOsP2jC3du0f3/GxWo1us7v+AxWW1
UhGYZy+mo903GpSd73+BHo1e9cS233pe/fta/aVhi9uK/7O7M2dS7ydAG3OfBt2A
CvX8dbbCDka7a+q3MiML5Pmkv7o9T6ETNYvMk+ankjcROL9Oc27A5m/LPxVhNLi8
D8DXD1H2W8BbfT68pGZwTRvDNas5/ZnYIe5VtZymWTNcVWgzaj5zl8cFBLYiYbv8
980ztwRDdclQPNNRk5QD1i9k9Gnlwv7p+z0RGVP1GgQqqv03DVNYnEg1lEDl4F2K
gdRj8pa9kmCmqFpB9EHVyqxWFD9WzLteQvkob/+sJzh7FTM5B9srfkkrjaUK+MH+
zLtmYgoKVjrTwhYjDFqMHoYk1WHrcmwbFEgzq43f+n3cKRBRK8UjAa9MR1mrsV5I
c1SPKRQB4vkPMDRYWKSGqS3S02AgQUcet2b5kbKRo7NcaQc/afiDbx2+v8utuCGQ
cTXRpzIO+u9JWyqYAope46W4ykf4Dbwd9u9fr8rkwozIx5TaihLKzMl0ZkExnLyt
DodyIAUlvX50uuurIQAqeaFE/IGBlRZkIOJmNwP6XdcpW8XAvRI2nx3WjH6o7F7H
YOPAtzP9X6pg8NlEOTkURjI4bxxUHKI2EDGRMJ5Va98T4qxbf9nIltP7f/9qPi7d
lbJPqdvQkyL/juNYzUUwQGfLmP8IXK5xtw05j0e8K35cKb2NZSBpIZ8OFRVMWcO1
SqXIEGNsIUqwhWexfb692Dskt3hEWDw8JaoIa4Juz5AksxpooKFan3s+3kTJWBNf
kev8AZGqdcfmIJHZJf0N2Ksy3IGeeAPeKbhjnfCQzXvIvHdFqtihI4iNknZjQOTG
O5tmLI6Qn7eOYE+3gGaoLJkhcQzi8EfxTwwLFOdpdItpS1QtJsti76xoQ3t59Cb0
o/gPZdtwFy3aNvVZBEJuJBROd8mk1VLoiVfgLp88E957x3latBptevfLtbD6RXxv
MZVmvx6G4TQBLANG81h5o8MeAktEekvU3EdD+7PArzakOyTgHmbM8AxT5KsMN4zg
34yVrOs2T7pjq9PZQeWzYmzsY1QNOHsljyISWUICaqaO1/CgLlfIc8B+0vxdfaSi
7Z8bBaAs4xSAwgWF3VOMha07IFb68Q2sokf4VJ/hf8tlbifCFozXqBjPml3ENlfT
6dTuJktW2tRijihxhPSewijE4TqLC9eX4vr2LsXymG0Ct0ZLOY1usVDCwIF3MA0B
jPTxHUVO5vgdhpxJRGFOiaph7+SkyNyZVN5p52BhOuPX/C15GkK/FhVjdqtQHkDN
AfW0jjJXWM15cNJqyKtoxllzK3+eMxzP4zULh6ntIT4i6JGPGbHo5KLhIAMLsRSH
7KPlUW0ODOBiNMICCiRF3n9j7s5CuxBDQdPZ2e2PhiYS9vq1AaiuT6q4srFmvmLv
LXgQFKMB+y8hJvmW3ufGCNtIGODS6i0ab2O8QIpvcDyz6QEGl4J90yDFZF5F1q99
nOgxeAexkYK9Urs6CoKW3xNAj6NMzV5e/J8M+Ez7ShEJykvub/uY6XUJtTh0errh
+bIqkXyJwlZXE4i44bxHeB/MnLPJAN/Gp29mzXqEE1e1afwj3ISNRCCkYh08+DYI
cNNAshhYs+kw1MJSx7grNU8rUdOeZNlNLclt/Zin6iFW3KtY34Bfq3O3rkY9gxSw
sb5hd8SujxdsnK4TGvuMEnlU5Rx3zSXsBkvimNZB8hA/O+xctC+0QftXn8sJY7B4
ff5RnMDHmznlQ4Dh6K2WWRii1ydEWJyyTwE5i82/lM/9gS4SNJMqnnXYvLp8/VWO
HTrUKyK0d0juDkbi0AorohsHGjf0cRvqhJMWIQ/H5fR70kyh4xU5ZZHxMCUAxz22
Jp185Y4hTZgNK/hMQ+fiCLqKJs59olGBpSkkw9airvepKMtyVihTKf8s2T2qFcHQ
o9HFe2f6EgjdAtxUgbwQf9mzOGs0Y608oKz3iR1hQu8XCk2DDw6ghEWo/2VwzBQH
kcXA4HCV8Y6Ds2NEapqZ6/rY+hTiTUQv6sJKGJxK3LTy1IZZIlumibg2qtXfgi9p
sC3aKtbMQ16zPngGrH4an7UElId8VnV0mFF+9ZxiMQbYjCGgKfJQG3KXepjax32n
MubWPicpH0vKJuw5FmLpE8345uGp4qrqQ1Q5l4I5GOitb74gBlwS37vyw4etsys9
ICWxyQT6SBitM/9pN6yvickQWEX9D3ir4+2wjBH2cFashK2+mGx2v6ww5VftMReS
KhdlC9D//stzQAV0uMmf/TpTac+21A+F1K0x6Lvsq3f08Oh3K842Jpiro8YoXsr3
lAQt2Oncg0gjqUFVQSI1/ZALX917vlFT8SYMUli/8MTvi5sTMdfCPlvIxDrKbrJ3
tx5P0Fq5CaJR2WyWeWikfB45dNpK6M6g2rkrLbJi+sgdeFK2jBkVbwDdJHi4Vjjn
y4nMd4r/ZY1RNaZ8bsIznkryH7aM7GnjA+Be6+3+DbXBucEgyo2EGXK1J/8GXjHY
WoyjwFFMkddzr3u5G6g02Z0DVz255uoSdBmVC8rnWf0e6b8hHnz+gtd+wwHLFojm
RTNGmQ8GeTqal6bnZFMcEdY6mGHKkIMEhQ4QRYUUOzyTpoAabXSIaBB2BDWPtuI+
RipD9DgDjNXGzs90dxaeuUMq+lSNA9JcWJUMODn66unjDulZOSKYygvab+3+tFyh
ttBsBKMod+zq0JQnd2uRbcJ5cF02kbE+wwUhKi0aGQMMxX1mlcKGyBmYGamBd7xb
0V0OIsjpMgYVSHTf+VXxe3B9Ljn49AFaNODXBcEU5aJQsp5Ye43fxvrNlM2yD2aM
IEtMHLOqldBN/Gbdnuo1yRkun1e+bGuEuBwh4l8dfs4H7DnizjN9Ww1FZcVp51tx
EYS9ENkwqTD7oAHvV7ioeqEMw+Z0xVtKODvV5JO2xNQWNTY+l7eNEdbt5Kr5qAbq
E6LDO6OUWWUy+b+LThZjuAGpH3dSZrN1p2ph1tRU0jZEwsdyx+Vg7GGM13PHrl2d
tHnQylL5HjtrQl5oyefC5m1v+C7r7bTbtaqGFD6imNfAPFx2x3n4jovMJrtJ0LbR
gecgWKIBg7VLJGlkG3ih12Qo3qu7NwpUXkchTnHPZ9vE5NLZNhPTbGzTfuxJXtuS
Uqg+QYd52MS9M782q11lBsFIty93eVb9a7/kNJPIpBFBhEsrVuEOfUBz9S0131hs
3tDU9zdY1ADpX/G5+4d0yDqitKbY/HBl3++sAnS3xaoyr/yztdqJeakDVdfp7hMQ
gVyeJHCPnKksmVE5vuOxhMXyWLr0I6JFvG18z7Yeq0l8l00jyQZGX24qSUQN8Grk
9y5lLIS3zhQhLMo7LbcUeDFlq1LFI0Tqn6qd0vGG4GafKbAqrnkhw10BhDtkDExs
gy1pvLL1mYvI82p9NDk9LAYtxC616+VARL6cO2cU7+oV0t8+qeAjbO/aWvdUXc2F
kxDc/UwjpMIaYQK5BOUh2Qq7Qc7sv78iFqdwhLi5NHC+MTjSWhbgkIdITO5lTFhn
WF2DROJ/xXy9e+ucK1S20Z29/iFzzMUmwAm7PPmorLCPaphIQbjCeESNgasFD8AF
7XwFRKlXIYQTVsWrL4lk0eKxVsWWBZEJnc7TyNk9UtVc0xzKAXmzsV8rUjKvBVRb
r6iIICc6UV5H3jqWJsmHj2olGfR1q6qiccYMua0xwiGFd5pMhcHLi4BFkO0D1BTe
PfJe/SP87/20Iyzz4wXFFLC8Gkhr/1rHPe71Ip9eKq5CU8bLVk39J9++fnKp8UqS
r2zEDayaSHtZkRjnAFVbZXeyh+2nlIZI9M4DO4gWDRFBA1OVog0aWeBE44CZJcZB
9mPcbqGOHqEilHsI116bCYVd8ITdRuVX8EtKP2AnBVBu4ZeC+Riwo+ZNsN6yfI6n
PdAHbJtFwed3J4v3RldShioKAKxMarfJnOgQf1poFuxwlJhN8o117t3OOT4gcx5S
wm+G0lpnaoK23QtUphBnc5Ja2Zzr2hoZ+oreeH0PjJJghkDdUQ2t+/sIEIbwcZLM
L09mZJFyVv0N20oESmzmck5UlOjW8DqCjoCnzdUJEayNYVrxxdzuHfplOQx6zHrR
UC/c7R9UFNF2/AXJxVk8s+o2+6Z+iFtPQFQ2x8aFjvpYUI6Ktk3atMPaLNeyoXLf
e2hKlEeV4Ojz7AZSFfw/V3AgS3Okm5r9EKy3nj+6rCnABM9X7F54SxW+A2vrsZo7
zbQj1pPd4datblgptDzLv+qWMKQLW6xoSahhgApbQ3n4H06W/b4dCBH0SaMYBbrP
viyF6LLcA8wnWid38WXTf2JdJHvOodjsdM13D2/NAhbyMLmkOScskkg59PKn2Isl
llXdCu3Rv7WddgOxqPApOw+gVUrEEq10npaRysXCkUmf6uuW9QfEFsyRkVmwqS/S
P1bP4N779gMF2rvVh9mSj+x8dXcm5hniLSr0AbF3SPo/LM99Ivb0zxqk2dYJWSeW
vR6ooIn9tkhJw1y6DKCes++r1rKrIGSmJc2zGvFr58t+HiwDMxSDgN3sTgGAC0gb
UNRsyg/HaxKVcZysHnl/KGbh0oD8/p1Atc/j76H6icfyLmL9kesH1Tsvarn76/pB
lQACLKZ+vpNKIzNOZCL/YAjDWkpdAXDTfNLsnlaLzA+QQiYLQ01EWz7odXoJ7jtf
PSQrnfTI4S7FutYgtHxsZxcIoi75sZnAXoch3aI0i6iJLDprYVFZHuMc4oVnjKg5
FLfKrEkKw1ofmA3jR1SwCcXrv0mcPFbj/hQeZII38EO0FCFNGROauXIxA2o8EJDm
y+FTdoVQ3x74Jo/4KMOFTwgWq5QGlI+o9qzsO50laKDlEb7/unfQNv/QyQoa75hk
Ir4bJgdIIYiPmyF3tA8u2vEijq81vYV+a7oQOt4QGiNiQRJK78y7Cx+wUQ/obEE/
XYbdIsmgN5CUM/Mq65gDG22VxIZsMd1PK4rxM2Vs0LymcQ5B5d3d9wp9U+ZPMFGn
skBu4gIjqa6Osi/uI0zTSxZyrMDpHy1Q4o1pL5NapS48I2QEJG+6bRssOXZutIoI
qEtGX+nYh86HGZZTdU6uFn9VZmHbwAA4GmjOOGn0TQzQ7e1RLZl7hStZzDFdTJsa
/GnjsWXZSbd6uC2k0FCExotCo1zwcgK7Znf658kwR9s=
`pragma protect end_protected
