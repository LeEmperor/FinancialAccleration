// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
G63Z1pUSXBVnX3wAA8UQbcrApux78k+uAE59mi6mi90ld2AgbTZL2G/XnlDRSFmutCQi2+zUFK41
qWGPQlR6nO/GeY8TGD5o8J0M8FCbvDUEEmnub45Qw58cX/V4biB54BXdQeViJ+/yY15THYt7AYUZ
JNR2EgzqSUWuHc3Q0LLbbbDwr7RJJZ1tSuw4gDnE26ZXz7tan6zM2Vyx4B1YVkF69rxAPlZ4BMGL
jzlFlbLuXpgHQaHV5yJvqRGsV962I+HNJdppFk7vJ8qSgGrjED6LuPB/lhp5obPdqc505dFiMj+j
frflBL1bDoTAEq90nXSOytODxkDCXkRRdV6HnQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
rpOsPpRJOOS5MxHFYsDTDvgXkRUnJyYUBUo7j2K6UgHib1ZjFesxmWND9W75cyH1ybXlB5fIoyoH
434XtCEMV0lslPiUn3RgICFX21vYrwf5aF3N9USFl8Z/Fl2LxqiqOUTbSh2FhgZUiqNFG7EzFb+D
wtBZS/wb5MEMwArmsFax1XPCULq6BR/EJWcoPFqZtqOT/KtFlRdMqH6iQAVQDwx5M9eO5bznTbjm
gzAhQVD+kxGH5+/FWrRjVUdhZVza9UwuPMV2iSSsQ8WnDr5PHuKmzyTkbtVWzSb837+l/ygTKVwY
aYfdB7Z22HzPc98wm31qISxjRUTFo1VY0Tbxy9JbdabNpK0QXLZa7eQ3E8Xv8UKBrvb8r04YVFE7
zomc3U6q1Zeb9ae0k0sQrpWbOZ4wWmgSse47F6RlOzxzaV5X79k5vjBXzoA8Gc9bUposEm4+iOX1
5W/wwLBSLKl7xBPJYTzuATLDUjy8mspNJ/9AElsSapzMPodJGUVP+yFhFliOCaNfdNGetuObPBXD
hB1Ksm+39bPJ9fAphX9wB6VsKuUMvmdmdQ0sf9rYQatsXje7fqPHgBpWaw4zWRZ9NTzVDp+3LNAq
4T1u0/NDitEdEED1hFyM5xAua5owWpVQjHGa53b30vLyHQ+zr0wrTaHC+Wa5KQfh202OAnbS/WzL
2Eg+W1kB7Na0eX9ag55RpGfTLx+rK2GJQD6rA2CethMJrJ9HwkzT7GIT677sEr+HQ67Pabzv91ht
gGf3RV4z2HZYeB/hsKw0twlBtj3DVL0IGXKcHOZC1w0JogGxsqPx0F7WoFrGj8DzG98VuBYV2my7
149zFUUeZIzcnw1EIT0nVW2VDsdSQbJbeBHuHzM6XAv0gCa5L4NoG0zaoKsryWiKeukBkDtS+wk8
3EtXdJIsBGxCJZoyBCupuav8ie/jtWJe3L7bmP5Ed6HQj0nq5XD+Iea9rsVbzf4Q/DadelwLZJqQ
9XbbJJOeP7QBSHPaDPGkI1fjWrRvOLmww6DVpPUQiath7mh0Qu3rrFcM9GixTveaW1VsWCcHDjvR
38Qj24C++ONmV3HTLuSy40KXJRw3fl/+85su0dkC8XtUhxQm1S0da6teVhlcvZF5Y6q9Fjfnmrls
syMR1GSmTP3J98B7a4O4MpjIBE+3tk0e2wFH2oTLOLfoMDg6nVPNwSeyfRo3CtlAcl1c/GUjr8DC
T2rC9icczB9/ngpDHZxlzpaf+yFX6mhGUs1SCxcFMZt+81Sakxwm4wKksRETzNNJgldF3oXDEBUM
rhK7GUrq+oTTGexyxawshdpuwnXR3hJgRNdM2Q0ll8vkKU520EUOJyaBo33AKz0jfujl5AV19l6+
4DpUT/TZ3VCQOL2VN9i6z+xnJHb5Cz8lCxnGm5FP105p9/1I6TYdASrrk1cM/jODiR1RA+4ZVtdb
wYK3pIIrQv2VO5bzZDH+eRxZCwgFVKKoCXcEb9ii5Hw+Rg1HY9FA/8sLXVhSFn9voV8BXDETJR8w
qRBjk8XnZnOonZFYTdr8pMPmCbD4W50CIuuZyad6lBM+5vUfbZPyJPwb/04eflRBXp6jppwChBtC
UEyOdCiMzNxZPuyDS+kZYYm7hNMqc13DKavmdRkJsSbN1Jbu1Dtx4xntKBm07yNMBLcfUUiRD3yQ
kdnLJJ180f3ESj9H8iwVxeni9cjqo/hUKqH44p5dPX9uTtZWM0AZsmX1uVST2M/X74VCBIzfShuN
+jy53ItZkctYgjAP4uwnVINv8gmRSUXq6E+Y8t/Jda26+asZiRCJEaNhL19tt/hpunGH0wqhZZ/o
Ql4HUgB5OYQnzEqHd10U9tuO/s9kZI3yCXlNatURF2wRU8GqTpxzWCzOQjwPpc+QKdr81oS6pgKd
chKMD2fkyBy0ZinvcIHFf0Wq9cXbMzqOlVtFkqSUqOp2LUFl1L7MTeugsyXEEQ9rNguq8n1G0T7R
jTRV6OSAOVLCZXN73u8GYELuVJ7+7bocXuJHcnVloS5ZtWMgPPu+maW0TaQZbagx8DHRzhO5vjgb
fMj+pZxLzG2PjsE2DA+pk1hpdT/JF/7ki+osfHZ4wLHMC1Co723p0ifFwbpkedq6LT4YEK3Sevnr
SfMtg3JLZCJcuGiJI66VavXAnPQdWIicv2XY5DVqXm5HsYTKcM3f2UAAe2zheScJAutjoaawtR3M
7rcIApvPP1d3w0OkyJxrjHiP4HHLUiDSQ6wLMBZIgj2d5v+48/36IiWmEQ/o9Bn9nwYFa/IDqQZK
eDNUsZ7ZMwlq63s9igR1bXOaMNhn8PGL5Eia/gADpq547GvA/wwE48bOow0jjkjd3FyySLTzWrkf
3CQ+I8t8akgiBKCgYLxcl6hgL2Rw0o7GtzZgzZFrGGPwaGQdi83QUEsNmUAm6/v0gjfl5l0J1viQ
qVUazHMwZYzjdTQwaCWtr/U79rDpRElhfIGMf6ZPhd9oGX7IPi2F2YAkXVWhQhttsJLkKB5EaRlo
wEdhvptKjpxBUDlZScIIMt43+DqmacMqkvXEQd6slrE7FSWw+eqD+z2zYNP13EhapEZEx16VwYLX
WpQIG7CmzQl7Y3anlw2qsJ6j5O/bUbA7dkaIZdawZViW64jD7gFQjaOCzkaLNg1HMXAxNESpWsoP
GRuZ5rVcAxA5tLKPrScmMMsZDkfNr3MW4RBbqOHZPfRN0QMOetpzebHeZpLLfb9sOfiQXVJdsViH
0+qAIH5oaSBOE7+K9MU92L4QmS/RN4hPv1m1sUmh9MyPkrooU0v/Qhz6IG1ZGb1YXKn/YoTpuzFo
KgErQUIyKAx3Y5+mfUqPZFNKeVD7JY43KcLZz2JgwpqfyISZzgGxfZpU+oHgeu7PdpSNYjYd2C6g
bjx/fVKYbxo4qags3nFFXKCYJhoxebR1Iex6vIU4u797Lkd0yI8Uhz2ArdxwdwqPbCYAGKoQM/8u
wbWH8P9KV49TXlivU6Ef+JmoJO1oka7No5fbdEGtPWgaow2sVSBCF/7OmqcbEJiuudZsmdWtHdBj
dFxFJu8ywQGUrrNgJavj7rEERE7MZuuFXlTgJZnOAZZV69QUrjQclNHimBGtPmTqAKWpfqTPGl8E
yST5WQv4wfByX1o+Et8/zK9WCV9XVJASDoRn4JaTtBEJXCPDEgUSOM0akIp3GWTDG77DEXh4ZgTQ
7zYMlUVRMaRtwhpC5Ay6vgBKqca0+emzcwqDgfAgDzcqyS5vGFitRNPum9S9UPhK/0fmGI5RvuWv
7ShEO2eDtH5H+muw8iFnyPTZp1ggtOlbeSop07C371Ix5hfzLEXdK/gMnVcu0Wd94bpQMXi1JJ/c
hdLLo0MTyfhUtWYo6oGKWbn6g3gMHthUXevMfeyKlyrdsilLum+UxSS1M9UU6MlDS4N0q0O/bWQE
RAxJhg/DnqqHCdHhozwDPT71SKDtIn6B+DKrpNAiLusrV2vKLWNTuDWJ7WPtZ8gDOGEs8VY6pwaB
CgB0GztC1y1IsnY+ecsU0VsBPSmZx0JsWuwR6sRc3K3ugmywLJQ+/vRS5h7xZcZ3bqusVPPIJ9XW
HzYgvKXZzBEWrrXyfM/HU0eo0e0LNFaz9YZv7Qkd8qGJQQH0aQuV3HYC3YWa0ZOgLhx4YOjP22qu
shyLoIKXcd2ZAYHFkiGKjpy2iZ1DMRUvg3CpjD7mcsl0hWPXX4R/OU2yNnYtu66liE4UWHp4b+xi
WQXoIJcj39vD9HSeHvVM6TGSa6+xYZuvWf9/W+cfWRHkGN1z0SRnynhXEOHUTkthv+7M/3YHKtws
EskSTB+rZrYlFQ2SPNn2XvhosBbYAvCtdO7uzS6rblb3zzDTR8LCDLbP70KeU8+nlVY8WLyRmL9n
QET5XQdNMossjQTxUa7/WMQrKldF321zCmWTpqaQpeHrbYMtRSdEriUHou4/cdL6BEIzZ8t9ZrYz
XBlrRk1drOffJ392nZbuLQN2EaDXUAj4rZThUQUv6fcGC8VQO3C2lNs3RWKNNCq8m/8m7nSJKpaR
v4tfgOyF1NIXvfNFx9R61BLugfJ2KOkwz0ZW8HVg5IiAr/1qC25FrpDEpAJMreOZTN/LDjbfWCi8
HB7Ugn0I5amZnRUonECBogJniCbjQfhgsWE9NVfX9ofpIEdc01vmu+ebQRz9DzmbDmDXA0OW4RyG
WaVZH8tG3VbYU+thoq1dyP6P2DH0FGpOG09m0mKt8QfucScVIbNr1dxVq/4F096yGjQI+Ef4vHDX
mgq+lChPrJL51SoZhblXpqahUuqAfgjNhxuFhdu6ESj6pyo5YAB62Ejqh69vsNcGr/v+IxrufnIM
DM0bHvnchdRMtUtqnabaTBw/a3LCelJSA/RDVjzMwauoFoi1B3+VrGNsL4FRKBOVEOlb1f8oQ75/
YznPbR+zNpahxjcfte64bYhilOvzRmPJUvp1WxfFCR0mD763NkKWKJA7wZCHgfTyizCUXF16MYJC
9GvlfRdLgvFpD5Fqi2103+m38cqsY6Dim6/2bl3gzORJv4YfC7hcZ7NmyM67GpdUj6V5HxJZlZGQ
gFJ3F9sfkQjOslF9F66kkKjZjT786xHKDo2UC4GMy9zOvmjb4Ua3M8OCqgimWeznTTZhKE/EVFqI
CVqQpckE9wWT75CQwc2HiXzR0g6FCa0FtYZ/y20nTrgYCa6mggsh7Tzr9MNiJe/jWWxvxIFmpJN4
mfcCIWj7BHmrK5pPg1XvqBfK1lwSQycH5aogGs66YBUAc1mp9tUgSK6cQtP6TpnJHry71tWMCcR5
KYprdRT7XeIvkFSQz3v9VCdYaRFCksrqz3I91fXLaYgCIuWVPQPFv779jtIjJcfRvBXoVg0JlmiK
4XdWQjs/83BkzsSaBah+GEpE8CAODPSTuCAmbb1mbyeP5lA2bdRHUuShpyuDcG4RZW/tw74/MuBc
jDqXgFu+37mfCbKKiaD7pDUif1AdykCBWTHO8yUkTRav5VG5T5QM6OyteSK+HUqTMdt7hSyS7mI6
1czqkzalAPUxl4+HwEin0MHU6MtoaRwAGUkebvUnZ/dduVU/1E1MgyMjv8FIoxJmukoJdGPc/6mS
3a4MsqEJhnI3dH7Qp1MhNN1xalEDSScT2bGSrOgVNAIO058wc/EpthAMve1d84UOPoSjXOVmCPeq
GXUZGK5Jy5vOsSwJ6eaZyNAtslu/sh1kD4n5g4l9iOOK+sv1nPqdjnK5+LbxKfN0Ah1JA9p9FwR8
R+iRrvCdoZeqMDGEzjfVHJJ+ibrXiz48MWBPr4qBdbglst8iJxy9y/H+OS2Wcr1NxFKVTvbQmSfM
75BztOgBbwXLYN1O1ONr0JtlKL2mAKFep3sdGMSV0qSuDAkBR9JURULUcCLBeEQO6BOmLpjKOzSQ
zqSlvzVk86BMfQMLmGjGXkeYyl/wD+awKmVcxPG3E/RwGP+Nj1B/85sEYtJA2MF1CmyjhzZ75L/J
HufaE5M5w03nlchvaONvDabwTwz1YFzX0TyHUVjeju9uuDmMeV98Xxw0fwYm0n+eXn+v+2rrQT52
dwUg87wu8IjnQug2cMXcimjy38i1zs3kolcmc52UPokZqS1r3BxSyoR3bJbmU8a+b2WqjSvypzt2
spvwrPY1D7aCQGRoRht5dN1MDgmlXTh+8odJkwpqsClCfKZ2XPm2qXipmuqG7OjjAWxN8WCcyXoB
wbbM+NP8yjkwu2H75u1YQ4pQCNZ0m++o8NNfocEbdC4AlCBa2ERD8PDE35tRAGE4o4HQREdlFZrG
+xT/nuEUfQ5j2liWVBcLkTZSIl4YXNSf7qo7XReNe90gsMCxh6KyETE387Hjw0v4hYA/V9gxlepb
UzjMetadMJF6yq4fNFXKZlzSQBJrlZOrLQnrNs0dRT4zn6INwOpzbWGKPJUKw0izTrr7Re6+MAc9
MRuH7LcjFB79rKaCj7YQb+Tm+Z1Pv7v7gam1U0d96uQsi6Gz0yGOSPLCf1xPOcAy47mvLrECupnh
yb7IQGQgDYe78bWgEIziJDKJ0m0OR/NoaNOq4ameXPObUNPL5I3oY04odvenkikuOrq3DHbOsUzE
zr9MyWdGGQPvvYqH9Z/yUUQSma8TMcq4x5hHdNF+A/DXFbilJy4vqOGhOvLLnEd4KdzCrKhIRaut
INC38mKzTtExNjLY6QV7R6yCDOX+/cGOkJ4bPAFI+eR6wmIpnQq2v/vp8SbT9Xu7hr0tYnCe4g94
imtjvY5l9fgdD5rB0YJmUIKGvq1Aec5wt1+7srtYGUJKEm/xZ9SN1ZzVa3gs+iKPLaD8GmaOQKe2
gQ6R3UDRor+te7ohKyBeSzSvCG31IC709wZDiHPAhzRZ9HDjZyUqMMT/SpNRd1sXDQ0FcFWeGKfq
5zuJnJhQoEY3xBWVLyn87qY7ugDZTgJb/HCiUdX1mT42gOH8XU0bKrtScm5bm0buDEcxXePvaF5b
lEiftOrSYc+nfvSoX3+H6cytba2S8AfJ4SQ5JLX0MYnpVZGZXlvizl459d8mdiK4vWeruLP4/MCe
afm2EAGac5QYUyzxLAEYQ/yaS9tjAKIhexOLzOJKv5slzKTBZ7VLUk7p/Af2IP71w0VNKOygBk/v
8ATKd0i3dlW1jZUqkuHL0Lq+iVau4n514MQIMkfYOLvb0otH04NbKFWgcPSTg2yOpkNKiG94FzY8
BmqknfCu+dix8l9vp4DE+tR+rDbtIIbr6nwN1Tt8rj9tYvZAW55jUFBYfhqEWr7DN3mBXy0W0Kr8
CDv9WcgT+H6BAGTqLZQBO7AL0yvTzI+jCWh72emnHwn2AzOVKDAbyu60r2Mh3L2QY1sK9x+YF4dU
jqJUJjdu5f54fdyez7g2NMmLaKRELPFJUIHMsLvFnTCynL98TCB+rA31MBlKgenuAIDA2bi80Byl
+MJdyTiM/iYFo0ihgzfWtmnyv8qW8xgUMny40uNAulvcUBFIfC5rvnB8QmnmYIRwozTH6FJwcrWb
8DYBOFpWFpZk1ndzZdMOB6q35ek=
`pragma protect end_protected
