`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CEntt2i0w1cXdKqw1RQUBj46k/U/HKimNSsIPkO0Hwvmma7Za3JjerRLm8XyIHiS
r4WmL/P3zE5+Xzu1FPUZG1Kn+6NAn89dfiBbNf+9IJUC/gPNMT2E8FGsZ4KL7pRd
I1v/mVtyuRitXx4RuIsQB1547hmQNpzxN2/58RAzgu0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
dKOghIUJMviK58X0pSkOLgpu84hzg3JTONlBnJLFRPZoNW6oxOseh8d1fsnX1ulJ
+HdSMirVmYZt8veGJ/3Sh0IGIhqGAavCfAsHnxHSEByDw0cEDfio9cB/OyGkOfmZ
Sg6yAg1o/ryprZqp7xpHNszN+MHJGuba4OdcdoLoAIqObIjqUZVdlHSMZup2VbIa
zY1Tvxu9Mz3pNNPQ2zsokGdBYGi2YrB59Yy7d2cMpKXQSjlA91qlSGqdlXxvVdP9
QIrOW+Jdka0pEJFBlZTIwvy1WJpVRCOaiR5sLz6vQq7XqpZCbkTr5yCEIWSqLn20
Oh4hlEV59prZvBRdULvFx7eHNmKfb2ZQjKKHwJiqp9qpQ8aNYZ0gxgsdHp6me0P2
YaK2p7ks4nuFioFz2j3i1ZDC7dqO/qc2NWE7OVAkfbRjvRtG6URijhzOYYkbpU7i
4/LwvanPd+OjX89WAHSD84dqyE19Wh9xyz6j2GPETfFthXxsteXcujaUpY4c/nG3
ODOl+3CXWLgbNyycIr/a4zWHXqPW5WwvZzPKU4YUowgYkryOlfXbii676PRjrXTt
UQioga2wW4AWkK6jlPfDlK6AT0O2PfNRw1xiu49UCtE9Or94jMZqTG1sQIAKfALH
dVN/+rjxJOmz7FYiT7ao2TFxhFTB2k7R2yZlQgH7fw5Huwi3hwdfeibtswHhFfbC
b+uzxbiPbTJ7Qy/aQMndOM3zmwdvZ8brjXEzEGCL7MXBtepe/0oPCNRvP/2lcn2h
e0jzIog8N1clyZU/ajm9/wlsEu0rUYSvZ6hwMNyOK07gTZyzDhY2tOEH2vJXmL/Y
E0uy5e0AEsEZUlLGVqSHuM7C+7cYSjV9EJF+pf1ESH+7+3n0b4CogRivySFUUVb4
l7d40odxaMABA0qp8dP4CHlU1NMSF31UflzKQW9Ry1dDjpOp2bS0OlUcf0c0w1Fa
bOZR4o2bFF29twYQOhITy6HwPO55UT6lnta3pwxyZewXVhH4yx+dQ5N1iRn8UxbY
oGgbSsVSp6XQ3ar8wbyI7LlaHECYLBAMVqst0bPbyyct629YIxEjfLYlrnA0qUX+
obY6I51+aQ1lkDI9KY5rtQtoYhcPmFZilFLGehowLX24/DwS3N4QVDkYxPJZGX0b
CnEFoO4FCZ+bwu4okROttDoeDDy/ZmGhjZiH7/K+NFoGthcSW2yvxjmzOobcwKp5
JSS8jntwPu/fakESye2mwgInLuTFQDxm2ATDhZc8Gv+k1eOoRltYnQLXWH4IHucv
r1/WweEZKJho35ShVwbMese3ncWx+d5fETIirzrcXmTkWdJq/jtl6h1r1xqJD3so
dYOe+0ypVTWWqKOXcPNV/45eS/5opKSqGB7h/p9aQHSKHPnO0MMqtJewoVznimv4
BNp/TK36ST41Dfacujeud2iFWyDldhVFFsfyqxlLbYZKs97TiybDVkdGeX5bTPjg
q2cnGNsOt2o34H9U+x9ZZ/H6VmlNp474H2YTnVs73xo3ib4UJSkL48jd9nC8dH6U
/VMZf75t/tHJi9bIrNosqsuqjuePOElywuY+79b4ctRxTuV1ETi65Iy78ARLqOI5
Itkt1oue1B2wS6+LLHWHr3nCIJTd0DNFEstJk0yyd6obP5rK4vQJy7Dp17X9Z8Mp
4JrR7JXOX+zuGVmgvCFzjdRflp47oTaEj50ZI9FNvKUuvd7uZ0+iYH7raYrSfJ/8
zOeswqFgJ3mhzgPEm+bAyGAn/J8az808X0m8RMaiOO50uO/mHbALBMlHCto7HyY5
gP3Et+3cJT0MEkFZyCF2JN3V2y9sFSquKzudMBcVkQQqbu8i/msKzXrBRMxMhFDF
OtpGLGq6A7FMRtHrUsa5PuUGSKIHdCHdQe2SFSvRLBS50TW1zO0EohDp98zRMLGL
IjbNE8ulfUYscZVufH4723B2H9c6mBAk3WQkpzIoRVqwp8sO8OZrpuANkl5UtQ0M
QcUjWHxYtsguzbfRD6RXkqcyjivz5uO+T+m9iQBwENxhkmN3gupGVeLqA/9EiD8b
f9loo2Nqb4VhhTjcBAq+khzuQ9tQg0x7/1sA4lMcyOgpnbCULF1FwVCBCjTvpih1
jUr6dx5ky5AwLNgzo+Fb34nkFs//D7uTR7mE8Fp2QupcuG+fzs4aiMfzOOWaRsAZ
dWE1ZMElZN4EBl7fsU3NpU4lgjEH5q2OIjuuqGK/XDpNgoO+f490D+zgxMRda/Ey
y20qV5Wvd3hJSU/bo9r+36k+Vjl7XpoRu1CsD6Tka8NvRb+Cu2FdET6bWiUkQWHX
MDch63rtOC5Cc+jo5/ixzUXgHYLfrd0tuLPhgyIHyvk0tU6gxVinVO6iZ/gj0BV1
abHrK58yLfbEX9Rp8jgGmzO2HuIPCbwLHFaZtTV0MfljTaCQquBRtJHtL3R68TsC
8yO4Nj0+ykX/jJxRfNyG42N0JsWAIeQ7shygU5SOdRpQu/nujtUNlnZ+87Vhs2qf
lM3VHf1gc/lAZFyi6wPcR1UBOmM1zcC1uKQLKw6bYQhA48EVCzfnPSqtwq3k9weg
gr8b5y/maJHH37VmL9y44AYVkYcK7uaDEKEbx7pjvDfliJErHh++UwSrMXhXajQ7
rvgk6c44QzueBM+6tvZIDFS/WIZ1XPQm9cn+LJZjp0cyN5Xseht4TeSzod1zjSn2
2BaTQlwPuuXf8rmNFfCjwp7ck6ET54ftiquzZgGGiubyb/i8qMmZfFJuOwQvHgdB
lwLHAmIkXntvX8kCYLZfBUZ6eAtIPUiPSH0WtcMy8B1CoREv2xx/+i/BnMQnPfKr
2EUVwyzbtMGQNGeirM5L9a57juJNRQYB2jRIax0/w4dbzhvJXuXUrp6P7eSkK0d/
+i6qD5eX+Kxyi+QXW4L9nHEfY+Xw1fRhMuxeCGPpPrVwB70wT2Qx0Et+ibcOGtLs
9hPCD9m5pWg8+tpEzN/IZweW02U1VvpJYx97xijZe676y41CVdPIoyj0CzIfewzL
g5mTlYtDfCT4dlmbkjKdGpfT0QxHhkN1BJXZi1jaaLqrVjaV0PyxDncRiJldussd
VK4p9jEn/iuWF//uEl9ad/ZtZtTQN7tt8FGgEpGUHzUCX/ZV/3+PRWd+AoYvv1/5
5VrLKpljdLB7TZ/2Zcl3SBxANY0jbauhtoI+XQ1MR7jJSIdd4xl1ahSVb6SDbSMH
dJwiK3katFycW3iV1Ih6SveujuX7WeuROw3B4F78Z3EZUxRuP0AVJZSfZy5k4ZRt
lFfrbzkcHDoNymZjjBnbL2I7Rp94LsJfePC4w5jr1gVgr61ELfLw0XLP0y5mlXN+
P2Xf/WAExpmIFEq7MLmMrCcoNkiH/2eDm3ZA/7sxBR3o7LaMt9xAxN50qOn4CCRA
Ba9OLsyqSIsqzXcRopcKe3wb/WdXWs4mlZKhQPd7rtZuzPZf7iOcBHfIs9QqJtIo
iZkUzWiXJKylr6preq6ufCpTXfo48F9MtnFrnvFQllELb8xzNEWkAlZRdnQdhzLy
P0eQObFKujS+FVboWx8Gfpjfn0xP4WjDuKRmHfUfV7rE2MAcbI0Q+ggujNkViUpG
H5eib93W1IY5UiuQ1AZnKRz/q67BcN/ksXcqKdcNqYcPt0gQboci2tk+D06FSbbm
uK9EERXGMhDuqQr14uoSRLazlxPGk5y69Xy4jB8eQpYuTziDHkFBS5DhTERg16Cy
MuAZa/ts04tVqnd2N4bDgMhsIRmyOK3SpQvkq8U8ws97IRFrpnae8spOTrS8NY/4
o3Sf8RnLEKgvv+Q7SvuburI3r4ByGf9oQq7tM4nFjS5rn6ma+/WIiMqSCrIxR+kR
XQrur3Bdo7YKV/zmcu9PLGODviKy4xntOBmptNzCLHOOcOcHhGGxIgkg1mu6xFxy
rDCocUlxz/GO1uQLGHxeFg35Asr9T7iy/kYMAr63ElsZEG2OxU8PEtNutUsbfO7M
aoiKNwjGRQJ3d+tSXx5PrMHtNF7VTB+NkUNa3Xr6EIG7TfACDE/1XScYiAhRtnim
h6+KRQceXOadzbOMKBr3S3Qe+If+gb2aWu7pwqvXR+KLWIFcZJJ8T3az782Ou7P+
RdVu7ZLRwR0KoJvzjSBFS46iT3r8F/VcAtQJNFwIdFzjOyzjP1Zgn+ryfdQ3MteX
JNfY6AKZ1FRSLEgOmmfcYMXjYenv6wF2axU+RvumGNHR5jIO2fpndSwhpSg36H5J
Kyr3E0XG2DXC9QjilncrmLyINxT55KZb5RKwbljpyX7dVyWT0ZEkOgD4gC+hhbqe
NXrbNi/PolyblQQu58nHmOa5JHU13NMCzPSDyEo+RIv7xKxBhbS18OaDy2K9sFsO
agXz2IG8QwUR1g4ixWRqtBxoaFOfKZV93Shp4x1+7a8L3UC7xeuWWv8V1WojsIoI
IaP2ijI9iYKkubSvDSZ32qLzGGdWOzOWksaQeZiGE81C1Skq/6PIk5hKn2UDrOuf
/oxX1kd89Jg5jPB1qyzl+lXloRDaIOf5G9GW2OydLkbWn87/RjEip9y2Zs62jWtL
77+UxE6oPr9m20N0wc7J696jvFFyXpmxn88gnMj0OHA1tCWhK4Sm0pZil/M0SRTb
LLFNS8sroT9ME97/XsYXCmlWQgZc8baJXKKtFGWFMdj6QfXbq2kiyYMtxIDPlDCB
QieA+8i+MvHGAlD9gnOlIwTVO+SMT84juxvEQIrqSmVGrUd0FFb2YMtLcnFs8CL5
i/4fX31ymAdPqPTj0AToU9TVCjhe1Ff0I3zNRQPaS4FxPF9nkZNeTNxX5G7tG8SX
hFfxTj9U6hW47q0D5AqbPzQzAP7QLR2FOlnZ6bCM6pbqtj5jcIc8ZeBC2y4SIQkw
boCjk9s9kqCybQjshsmDZsyYCtPS4NxGB3sGZPW3JSbZBtAm10AupaZ8AlIBtQV/
GtkMATgXqNG4C6ECSl0rkDuZBovrtLUrD1CisK7iTl3cVWu9CGDEIxW1bhcmGnPG
CVjaU6YFYFqJ8DA+6KHzEMd5lC8qxGQuDz2lBPh0+GVncfiy0NP4pzXtXSvXn01f
lU+8hJ2pgVuS+Jh+hMm/LtAUVI/91PSJcAXPrMiZYln1jQP5s2MBR8gIbABBE/59
mrx65AdYoumGWkBn0v/nf1CcrGSpzRUFP28lLh54qsh2suSmwJGnScCVkPQ0WmUO
wj+E0ouAc0J4CyxRRGc2/+isRSkBKA+XCm+u38tqQXbirlt4lAcbrsRNrICgfDHr
g//yVKsjtSBK/MU0tKOHyhBAMwoHl4tMt2Ve6amCmYD5uHVnKACuiW7JRrQ+B8tt
go/NDpvOeC/xdPOfVoWom0PEdMXqgrA1Qk/Tfh68EKiPbwGKT2v7wi82XwbKfZBk
wZCTWYh5fiWrMKRUBETkdsJqrUflXg0/zyoCBDCepCXQVICyRe2IS8GT3Z4r7dAe
vmvE0nNo30r4D0nqaoU3rwAAjxTWt3IVXqw1SIr9OGPLAcr/l0jzG6tQsdjssonu
OvMKa2EmMVPsVN8qAHV0Xt2zWMLThpy/NhLNlN8Vyfe90cWUvWu6VkeRWJ0DmmFB
JNUQ/XmLWAAdNLcSUzLo1NeT/7uGRCe8ArIjPoEBlFwcxdsOVqQ/EzhB/dwoHQIy
SlBjJaOiQ5QpiEJPpMD9UIB8Sf5P+yYqy8RIMpc8/7ujDf8Le1uQ7cy1G1s770sG
r8UJorP6ZdbTyXOTLz03gHkMw7xaVA6/7KzsjCA2DHZNHQl6ezl1rQSAqtFf61pW
lGjDzlzGETC5wZaoQOvkFkJbmBXyNG8MRyKM15OGQ9uMpo7ot2hk0YNNifOWRjGI
T3fEKrpE7t6j2RzMnUPHP7mwE8civl0dwu/CcGlQM/rggxzfJ8VKYni5CcZSRGI1
9Tlks5kqh8RHhOt4C5DzpeI10TLdHQ9dK+P4Xshxbaejl7AirZ0TMQfkYU4/QQHf
dRAYgG760TbEpR+njzlbMnvZyJwk7o2lJ/xa9VB7x6eXSy+EvBusr+CI+35LLv7p
k46HMmR6caEGeW1IqFz13wVkMk71nausBpVhMgEdyJSZcTavVbgczfELWJm8ks59
jB5Dp/uWyyU5Xug3M8n9iGKCDAH1d0BzyDFRnwdyzzrYfmG4V2h10ehrdxUclnoe
7DnhTOlv1sW8HHlNVTAV4ZJxtJDTtsKP6wjth/KTa8GHaSnlD7g9SI9ShwAhtptV
5zk7VhTSgz1ajqkCWYgLXf8HsubEOrzFnc4U+kyP+mtYwzhvwiPwrBAYxb/mWi3f
MjmX6ji6lDNJ/itKbLZgZsanhmBadc4o3lsKFCJm7pMxm2kTUby3uQfy8Q0plkB9
nAouzS7TzGALC13frKFcvieVKe35wnxd1wfwzS/MllKMPK94B6HXE503LTfbnYLn
5mREZYM2IFEvvsIzGj2DzORiEc3KaSv33mSG8R4pi5r6TiiOoi1KZ/xrPxBAn23R
tdiLR7nwaak+ht9flgJ4XQ3l+j2KE/r+XialKjI8nEdL5AVGZCHdtF7BSUSc4gJ2
2x3NnInHY3dAjfkaybHFVj2xrsYNCPxkcejYc8VSADcSop1nwlzs0tuRoljixFrq
Tgzc8Jr7xcmCAg7jKhQH3JIdKSvlNZF99aNwt8qItUn67jBn9n1tk1eJx8t2RLP9
Ni2CLYpZB/cqoEtlmu0vZjbUopMTcnkMv3zUJVGzAjBIt+jSmhAM+3gO9+p7l/JV
cf3QNxNMCCfc2ymtiamY1RzSBNbrXDv5wffMvrSIhFNW2ikL/g81uGD7qdX0Kdiu
ytRvzVEIPRPhAOW65z3QzHcVEPaVZ0XHVewuViYm9FGORDL00J6+A+gVls6IEv2f
NiRk+s6uBovrwYlXxxPMi4Zx6RcvmLAXCrnB37+uFC5ggQNHXHTuYwPTWDRCP0UV
3aICmcOVpzWs7BmLN++hJADkTovfn7BiNz6v2jQLImxgVJLC2TLtwI7LkMXqXbgM
OiGPUBJlkzL7pShhfJQwzf4MwmgIoaOFYwSaKQH+pymUJ3yqZUGs7n6m5SqDCYO6
+MZ10Fvf5NgkLPkl+2TC6BTlhoIBeKR/PKFIcbPJQC7DAEu4RXImSVKgvK7+JLti
59g3k4+l4ytSZqLYzIN3KA==
`pragma protect end_protected
